
module acc_user_1 #
(
  parameter DATA_WIDTH = 32,
  parameter NUM_INPUT_QUEUES = 1,
  parameter NUM_OUTPUT_QUEUES = 1
)
(
  input clk,
  input rst,
  input start,
  input [2-1:0] acc_user_done_rd_data,
  input [2-1:0] acc_user_done_wr_data,
  input [2-1:0] acc_user_available_read,
  input [1024-1:0] acc_user_read_data,
  output [2-1:0] acc_user_request_read,
  input [2-1:0] acc_user_read_data_valid,
  input [2-1:0] acc_user_available_write,
  output [1024-1:0] acc_user_write_data,
  output [2-1:0] acc_user_request_write,
  output reg acc_user_done
);

  wire [34-1:0] n0;
  wire [34-1:0] n1;
  wire [34-1:0] n10;
  wire [34-1:0] n100;
  wire [34-1:0] n1000;
  wire [34-1:0] n1001;
  wire [34-1:0] n1002;
  wire [34-1:0] n1003;
  wire [34-1:0] n1004;
  wire [34-1:0] n1005;
  wire [34-1:0] n1006;
  wire [34-1:0] n1007;
  wire [34-1:0] n1008;
  wire [34-1:0] n1009;
  wire [34-1:0] n101;
  wire [34-1:0] n1010;
  wire [34-1:0] n1011;
  wire [34-1:0] n1012;
  wire [34-1:0] n1013;
  wire [34-1:0] n1014;
  wire [34-1:0] n1015;
  wire [34-1:0] n1016;
  wire [34-1:0] n1017;
  wire [34-1:0] n1018;
  wire [34-1:0] n1019;
  wire [34-1:0] n102;
  wire [34-1:0] n1020;
  wire [34-1:0] n1021;
  wire [34-1:0] n1022;
  wire [34-1:0] n1023;
  wire [34-1:0] n1024;
  wire [34-1:0] n1025;
  wire [34-1:0] n1026;
  wire [34-1:0] n1027;
  wire [34-1:0] n1028;
  wire [34-1:0] n1029;
  wire [34-1:0] n103;
  wire [34-1:0] n1030;
  wire [34-1:0] n1031;
  wire [34-1:0] n1032;
  wire [34-1:0] n1033;
  wire [34-1:0] n1034;
  wire [34-1:0] n1035;
  wire [34-1:0] n1036;
  wire [34-1:0] n1037;
  wire [34-1:0] n1038;
  wire [34-1:0] n1039;
  wire [34-1:0] n104;
  wire [34-1:0] n1040;
  wire [34-1:0] n1041;
  wire [34-1:0] n1042;
  wire [34-1:0] n1043;
  wire [34-1:0] n1044;
  wire [34-1:0] n1045;
  wire [34-1:0] n1046;
  wire [34-1:0] n1047;
  wire [34-1:0] n1048;
  wire [34-1:0] n1049;
  wire [34-1:0] n105;
  wire [34-1:0] n1050;
  wire [34-1:0] n1051;
  wire [34-1:0] n1052;
  wire [34-1:0] n1053;
  wire [34-1:0] n1054;
  wire [34-1:0] n1055;
  wire [34-1:0] n1056;
  wire [34-1:0] n1057;
  wire [34-1:0] n1058;
  wire [34-1:0] n1059;
  wire [34-1:0] n106;
  wire [34-1:0] n1060;
  wire [34-1:0] n1061;
  wire [34-1:0] n1062;
  wire [34-1:0] n1063;
  wire [34-1:0] n1064;
  wire [34-1:0] n1065;
  wire [34-1:0] n1066;
  wire [34-1:0] n1067;
  wire [34-1:0] n1068;
  wire [34-1:0] n1069;
  wire [34-1:0] n107;
  wire [34-1:0] n1070;
  wire [34-1:0] n1071;
  wire [34-1:0] n1072;
  wire [34-1:0] n1073;
  wire [34-1:0] n1074;
  wire [34-1:0] n1075;
  wire [34-1:0] n1076;
  wire [34-1:0] n1077;
  wire [34-1:0] n1078;
  wire [34-1:0] n1079;
  wire [34-1:0] n108;
  wire [34-1:0] n1080;
  wire [34-1:0] n1081;
  wire [34-1:0] n1082;
  wire [34-1:0] n1083;
  wire [34-1:0] n1084;
  wire [34-1:0] n1085;
  wire [34-1:0] n1086;
  wire [34-1:0] n1087;
  wire [34-1:0] n1088;
  wire [34-1:0] n1089;
  wire [34-1:0] n109;
  wire [34-1:0] n1090;
  wire [34-1:0] n1091;
  wire [34-1:0] n1092;
  wire [34-1:0] n1093;
  wire [34-1:0] n1094;
  wire [34-1:0] n1095;
  wire [34-1:0] n1096;
  wire [34-1:0] n1097;
  wire [34-1:0] n1098;
  wire [34-1:0] n1099;
  wire [34-1:0] n11;
  wire [34-1:0] n110;
  wire [34-1:0] n1100;
  wire [34-1:0] n1101;
  wire [34-1:0] n1102;
  wire [34-1:0] n1103;
  wire [34-1:0] n1104;
  wire [34-1:0] n1105;
  wire [34-1:0] n1106;
  wire [34-1:0] n1107;
  wire [34-1:0] n1108;
  wire [34-1:0] n1109;
  wire [34-1:0] n111;
  wire [34-1:0] n1110;
  wire [34-1:0] n1111;
  wire [34-1:0] n1112;
  wire [34-1:0] n1113;
  wire [34-1:0] n1114;
  wire [34-1:0] n1115;
  wire [34-1:0] n1116;
  wire [34-1:0] n1117;
  wire [34-1:0] n1118;
  wire [34-1:0] n1119;
  wire [34-1:0] n112;
  wire [34-1:0] n1120;
  wire [34-1:0] n1121;
  wire [34-1:0] n1122;
  wire [34-1:0] n1123;
  wire [34-1:0] n1124;
  wire [34-1:0] n1125;
  wire [34-1:0] n1126;
  wire [34-1:0] n1127;
  wire [34-1:0] n1128;
  wire [34-1:0] n1129;
  wire [34-1:0] n113;
  wire [34-1:0] n1130;
  wire [34-1:0] n1131;
  wire [34-1:0] n1132;
  wire [34-1:0] n1133;
  wire [34-1:0] n1134;
  wire [34-1:0] n1135;
  wire [34-1:0] n1136;
  wire [34-1:0] n1137;
  wire [34-1:0] n1138;
  wire [34-1:0] n1139;
  wire [34-1:0] n114;
  wire [34-1:0] n1140;
  wire [34-1:0] n1141;
  wire [34-1:0] n1142;
  wire [34-1:0] n1143;
  wire [34-1:0] n1144;
  wire [34-1:0] n1145;
  wire [34-1:0] n1146;
  wire [34-1:0] n1147;
  wire [34-1:0] n1148;
  wire [34-1:0] n1149;
  wire [34-1:0] n115;
  wire [34-1:0] n1150;
  wire [34-1:0] n1151;
  wire [34-1:0] n1152;
  wire [34-1:0] n1153;
  wire [34-1:0] n1154;
  wire [34-1:0] n1155;
  wire [34-1:0] n1156;
  wire [34-1:0] n1157;
  wire [34-1:0] n1158;
  wire [34-1:0] n1159;
  wire [34-1:0] n116;
  wire [34-1:0] n1160;
  wire [34-1:0] n1161;
  wire [34-1:0] n1162;
  wire [34-1:0] n1163;
  wire [34-1:0] n1164;
  wire [34-1:0] n1165;
  wire [34-1:0] n1166;
  wire [34-1:0] n1167;
  wire [34-1:0] n1168;
  wire [34-1:0] n1169;
  wire [34-1:0] n117;
  wire [34-1:0] n1170;
  wire [34-1:0] n1171;
  wire [34-1:0] n1172;
  wire [34-1:0] n1173;
  wire [34-1:0] n1174;
  wire [34-1:0] n1175;
  wire [34-1:0] n1176;
  wire [34-1:0] n1177;
  wire [34-1:0] n1178;
  wire [34-1:0] n1179;
  wire [34-1:0] n118;
  wire [34-1:0] n1180;
  wire [34-1:0] n1181;
  wire [34-1:0] n1182;
  wire [34-1:0] n1183;
  wire [34-1:0] n1184;
  wire [34-1:0] n1185;
  wire [34-1:0] n1186;
  wire [34-1:0] n1187;
  wire [34-1:0] n1188;
  wire [34-1:0] n1189;
  wire [34-1:0] n119;
  wire [34-1:0] n1190;
  wire [34-1:0] n1191;
  wire [34-1:0] n1192;
  wire [34-1:0] n1193;
  wire [34-1:0] n1194;
  wire [34-1:0] n1195;
  wire [34-1:0] n1196;
  wire [34-1:0] n1197;
  wire [34-1:0] n1198;
  wire [34-1:0] n1199;
  wire [34-1:0] n12;
  wire [34-1:0] n120;
  wire [34-1:0] n1200;
  wire [34-1:0] n1201;
  wire [34-1:0] n1202;
  wire [34-1:0] n1203;
  wire [34-1:0] n1204;
  wire [34-1:0] n1205;
  wire [34-1:0] n1206;
  wire [34-1:0] n1207;
  wire [34-1:0] n1208;
  wire [34-1:0] n1209;
  wire [34-1:0] n121;
  wire [34-1:0] n1210;
  wire [34-1:0] n1211;
  wire [34-1:0] n1212;
  wire [34-1:0] n1213;
  wire [34-1:0] n1214;
  wire [34-1:0] n1215;
  wire [34-1:0] n1216;
  wire [34-1:0] n1217;
  wire [34-1:0] n1218;
  wire [34-1:0] n1219;
  wire [34-1:0] n122;
  wire [34-1:0] n1220;
  wire [34-1:0] n1221;
  wire [34-1:0] n1222;
  wire [34-1:0] n1223;
  wire [34-1:0] n1224;
  wire [34-1:0] n1225;
  wire [34-1:0] n1226;
  wire [34-1:0] n1227;
  wire [34-1:0] n1228;
  wire [34-1:0] n1229;
  wire [34-1:0] n123;
  wire [34-1:0] n1230;
  wire [34-1:0] n1231;
  wire [34-1:0] n1232;
  wire [34-1:0] n1233;
  wire [34-1:0] n1234;
  wire [34-1:0] n1235;
  wire [34-1:0] n1236;
  wire [34-1:0] n1237;
  wire [34-1:0] n1238;
  wire [34-1:0] n1239;
  wire [34-1:0] n124;
  wire [34-1:0] n1240;
  wire [34-1:0] n1241;
  wire [34-1:0] n1242;
  wire [34-1:0] n1243;
  wire [34-1:0] n1244;
  wire [34-1:0] n1245;
  wire [34-1:0] n1246;
  wire [34-1:0] n1247;
  wire [34-1:0] n1248;
  wire [34-1:0] n1249;
  wire [34-1:0] n125;
  wire [34-1:0] n1250;
  wire [34-1:0] n1251;
  wire [34-1:0] n1252;
  wire [34-1:0] n1253;
  wire [34-1:0] n1254;
  wire [34-1:0] n1255;
  wire [34-1:0] n1256;
  wire [34-1:0] n1257;
  wire [34-1:0] n1258;
  wire [34-1:0] n1259;
  wire [34-1:0] n126;
  wire [34-1:0] n1260;
  wire [34-1:0] n1261;
  wire [34-1:0] n1262;
  wire [34-1:0] n1263;
  wire [34-1:0] n1264;
  wire [34-1:0] n1265;
  wire [34-1:0] n1266;
  wire [34-1:0] n1267;
  wire [34-1:0] n1268;
  wire [34-1:0] n1269;
  wire [34-1:0] n127;
  wire [34-1:0] n1270;
  wire [34-1:0] n1271;
  wire [34-1:0] n1272;
  wire [34-1:0] n1273;
  wire [34-1:0] n1274;
  wire [34-1:0] n1275;
  wire [34-1:0] n1276;
  wire [34-1:0] n1277;
  wire [34-1:0] n1278;
  wire [34-1:0] n1279;
  wire [34-1:0] n128;
  wire [34-1:0] n1280;
  wire [34-1:0] n1281;
  wire [34-1:0] n1282;
  wire [34-1:0] n1283;
  wire [34-1:0] n1284;
  wire [34-1:0] n1285;
  wire [34-1:0] n1286;
  wire [34-1:0] n1287;
  wire [34-1:0] n1288;
  wire [34-1:0] n1289;
  wire [34-1:0] n129;
  wire [34-1:0] n1290;
  wire [34-1:0] n1291;
  wire [34-1:0] n1292;
  wire [34-1:0] n1293;
  wire [34-1:0] n1294;
  wire [34-1:0] n1295;
  wire [34-1:0] n1296;
  wire [34-1:0] n1297;
  wire [34-1:0] n1298;
  wire [34-1:0] n1299;
  wire [34-1:0] n13;
  wire [34-1:0] n130;
  wire [34-1:0] n1300;
  wire [34-1:0] n1301;
  wire [34-1:0] n1302;
  wire [34-1:0] n1303;
  wire [34-1:0] n1304;
  wire [34-1:0] n1305;
  wire [34-1:0] n1306;
  wire [34-1:0] n1307;
  wire [34-1:0] n1308;
  wire [34-1:0] n1309;
  wire [34-1:0] n131;
  wire [34-1:0] n1310;
  wire [34-1:0] n1311;
  wire [34-1:0] n1312;
  wire [34-1:0] n1313;
  wire [34-1:0] n1314;
  wire [34-1:0] n1315;
  wire [34-1:0] n1316;
  wire [34-1:0] n1317;
  wire [34-1:0] n1318;
  wire [34-1:0] n1319;
  wire [34-1:0] n132;
  wire [34-1:0] n1320;
  wire [34-1:0] n1321;
  wire [34-1:0] n1322;
  wire [34-1:0] n1323;
  wire [34-1:0] n1324;
  wire [34-1:0] n1325;
  wire [34-1:0] n1326;
  wire [34-1:0] n1327;
  wire [34-1:0] n1328;
  wire [34-1:0] n1329;
  wire [34-1:0] n133;
  wire [34-1:0] n1330;
  wire [34-1:0] n1331;
  wire [34-1:0] n1332;
  wire [34-1:0] n1333;
  wire [34-1:0] n1334;
  wire [34-1:0] n1335;
  wire [34-1:0] n1336;
  wire [34-1:0] n1337;
  wire [34-1:0] n1338;
  wire [34-1:0] n1339;
  wire [34-1:0] n134;
  wire [34-1:0] n1340;
  wire [34-1:0] n1341;
  wire [34-1:0] n1342;
  wire [34-1:0] n1343;
  wire [34-1:0] n1344;
  wire [34-1:0] n1345;
  wire [34-1:0] n1346;
  wire [34-1:0] n1347;
  wire [34-1:0] n1348;
  wire [34-1:0] n1349;
  wire [34-1:0] n135;
  wire [34-1:0] n1350;
  wire [34-1:0] n1351;
  wire [34-1:0] n1352;
  wire [34-1:0] n1353;
  wire [34-1:0] n1354;
  wire [34-1:0] n1355;
  wire [34-1:0] n1356;
  wire [34-1:0] n1357;
  wire [34-1:0] n1358;
  wire [34-1:0] n1359;
  wire [34-1:0] n136;
  wire [34-1:0] n1360;
  wire [34-1:0] n1361;
  wire [34-1:0] n1362;
  wire [34-1:0] n1363;
  wire [34-1:0] n1364;
  wire [34-1:0] n1365;
  wire [34-1:0] n1366;
  wire [34-1:0] n1367;
  wire [34-1:0] n1368;
  wire [34-1:0] n1369;
  wire [34-1:0] n137;
  wire [34-1:0] n1370;
  wire [34-1:0] n1371;
  wire [34-1:0] n1372;
  wire [34-1:0] n1373;
  wire [34-1:0] n1374;
  wire [34-1:0] n1375;
  wire [34-1:0] n1376;
  wire [34-1:0] n1377;
  wire [34-1:0] n1378;
  wire [34-1:0] n1379;
  wire [34-1:0] n138;
  wire [34-1:0] n1380;
  wire [34-1:0] n1381;
  wire [34-1:0] n1382;
  wire [34-1:0] n1383;
  wire [34-1:0] n1384;
  wire [34-1:0] n1385;
  wire [34-1:0] n1386;
  wire [34-1:0] n1387;
  wire [34-1:0] n1388;
  wire [34-1:0] n1389;
  wire [34-1:0] n139;
  wire [34-1:0] n1390;
  wire [34-1:0] n1391;
  wire [34-1:0] n1392;
  wire [34-1:0] n1393;
  wire [34-1:0] n1394;
  wire [34-1:0] n1395;
  wire [34-1:0] n1396;
  wire [34-1:0] n1397;
  wire [34-1:0] n1398;
  wire [34-1:0] n1399;
  wire [34-1:0] n14;
  wire [34-1:0] n140;
  wire [34-1:0] n1400;
  wire [34-1:0] n1401;
  wire [34-1:0] n1402;
  wire [34-1:0] n1403;
  wire [34-1:0] n1404;
  wire [34-1:0] n1405;
  wire [34-1:0] n1406;
  wire [34-1:0] n1407;
  wire [34-1:0] n1408;
  wire [34-1:0] n1409;
  wire [34-1:0] n141;
  wire [34-1:0] n1410;
  wire [34-1:0] n1411;
  wire [34-1:0] n1412;
  wire [34-1:0] n1413;
  wire [34-1:0] n1414;
  wire [34-1:0] n1415;
  wire [34-1:0] n1416;
  wire [34-1:0] n1417;
  wire [34-1:0] n1418;
  wire [34-1:0] n1419;
  wire [34-1:0] n142;
  wire [34-1:0] n1420;
  wire [34-1:0] n1421;
  wire [34-1:0] n1422;
  wire [34-1:0] n1423;
  wire [34-1:0] n1424;
  wire [34-1:0] n1425;
  wire [34-1:0] n1426;
  wire [34-1:0] n1427;
  wire [34-1:0] n1428;
  wire [34-1:0] n1429;
  wire [34-1:0] n143;
  wire [34-1:0] n1430;
  wire [34-1:0] n1431;
  wire [34-1:0] n1432;
  wire [34-1:0] n1433;
  wire [34-1:0] n1434;
  wire [34-1:0] n1435;
  wire [34-1:0] n1436;
  wire [34-1:0] n1437;
  wire [34-1:0] n1438;
  wire [34-1:0] n1439;
  wire [34-1:0] n144;
  wire [34-1:0] n1440;
  wire [34-1:0] n1441;
  wire [34-1:0] n1442;
  wire [34-1:0] n1443;
  wire [34-1:0] n1444;
  wire [34-1:0] n1445;
  wire [34-1:0] n1446;
  wire [34-1:0] n1447;
  wire [34-1:0] n1448;
  wire [34-1:0] n1449;
  wire [34-1:0] n145;
  wire [34-1:0] n1450;
  wire [34-1:0] n1451;
  wire [34-1:0] n1452;
  wire [34-1:0] n1453;
  wire [34-1:0] n1454;
  wire [34-1:0] n1455;
  wire [34-1:0] n1456;
  wire [34-1:0] n1457;
  wire [34-1:0] n1458;
  wire [34-1:0] n1459;
  wire [34-1:0] n146;
  wire [34-1:0] n1460;
  wire [34-1:0] n1461;
  wire [34-1:0] n1462;
  wire [34-1:0] n1463;
  wire [34-1:0] n1464;
  wire [34-1:0] n1465;
  wire [34-1:0] n1466;
  wire [34-1:0] n1467;
  wire [34-1:0] n1468;
  wire [34-1:0] n1469;
  wire [34-1:0] n147;
  wire [34-1:0] n1470;
  wire [34-1:0] n1471;
  wire [34-1:0] n1472;
  wire [34-1:0] n1473;
  wire [34-1:0] n1474;
  wire [34-1:0] n1475;
  wire [34-1:0] n1476;
  wire [34-1:0] n1477;
  wire [34-1:0] n1478;
  wire [34-1:0] n1479;
  wire [34-1:0] n148;
  wire [34-1:0] n1480;
  wire [34-1:0] n1481;
  wire [34-1:0] n1482;
  wire [34-1:0] n1483;
  wire [34-1:0] n1484;
  wire [34-1:0] n1485;
  wire [34-1:0] n1486;
  wire [34-1:0] n1487;
  wire [34-1:0] n1488;
  wire [34-1:0] n1489;
  wire [34-1:0] n149;
  wire [34-1:0] n1490;
  wire [34-1:0] n1491;
  wire [34-1:0] n1492;
  wire [34-1:0] n1493;
  wire [34-1:0] n1494;
  wire [34-1:0] n1495;
  wire [34-1:0] n1496;
  wire [34-1:0] n1497;
  wire [34-1:0] n1498;
  wire [34-1:0] n1499;
  wire [34-1:0] n15;
  wire [34-1:0] n150;
  wire [34-1:0] n1500;
  wire [34-1:0] n1501;
  wire [34-1:0] n1502;
  wire [34-1:0] n1503;
  wire [34-1:0] n1504;
  wire [34-1:0] n1505;
  wire [34-1:0] n1506;
  wire [34-1:0] n1507;
  wire [34-1:0] n1508;
  wire [34-1:0] n1509;
  wire [34-1:0] n151;
  wire [34-1:0] n1510;
  wire [34-1:0] n1511;
  wire [34-1:0] n1512;
  wire [34-1:0] n1513;
  wire [34-1:0] n1514;
  wire [34-1:0] n1515;
  wire [34-1:0] n1516;
  wire [34-1:0] n1517;
  wire [34-1:0] n1518;
  wire [34-1:0] n1519;
  wire [34-1:0] n152;
  wire [34-1:0] n1520;
  wire [34-1:0] n1521;
  wire [34-1:0] n1522;
  wire [34-1:0] n1523;
  wire [34-1:0] n1524;
  wire [34-1:0] n1525;
  wire [34-1:0] n1526;
  wire [34-1:0] n1527;
  wire [34-1:0] n1528;
  wire [34-1:0] n1529;
  wire [34-1:0] n153;
  wire [34-1:0] n1530;
  wire [34-1:0] n1531;
  wire [34-1:0] n1532;
  wire [34-1:0] n1533;
  wire [34-1:0] n1534;
  wire [34-1:0] n1535;
  wire [34-1:0] n1536;
  wire [34-1:0] n1537;
  wire [34-1:0] n1538;
  wire [34-1:0] n1539;
  wire [34-1:0] n154;
  wire [34-1:0] n1540;
  wire [34-1:0] n1541;
  wire [34-1:0] n1542;
  wire [34-1:0] n1543;
  wire [34-1:0] n1544;
  wire [34-1:0] n1545;
  wire [34-1:0] n1546;
  wire [34-1:0] n1547;
  wire [34-1:0] n1548;
  wire [34-1:0] n1549;
  wire [34-1:0] n155;
  wire [34-1:0] n1550;
  wire [34-1:0] n1551;
  wire [34-1:0] n1552;
  wire [34-1:0] n1553;
  wire [34-1:0] n1554;
  wire [34-1:0] n1555;
  wire [34-1:0] n1556;
  wire [34-1:0] n1557;
  wire [34-1:0] n1558;
  wire [34-1:0] n1559;
  wire [34-1:0] n156;
  wire [34-1:0] n1560;
  wire [34-1:0] n1561;
  wire [34-1:0] n1562;
  wire [34-1:0] n1563;
  wire [34-1:0] n1564;
  wire [34-1:0] n1565;
  wire [34-1:0] n1566;
  wire [34-1:0] n1567;
  wire [34-1:0] n1568;
  wire [34-1:0] n1569;
  wire [34-1:0] n157;
  wire [34-1:0] n1570;
  wire [34-1:0] n1571;
  wire [34-1:0] n1572;
  wire [34-1:0] n1573;
  wire [34-1:0] n1574;
  wire [34-1:0] n1575;
  wire [34-1:0] n1576;
  wire [34-1:0] n1577;
  wire [34-1:0] n1578;
  wire [34-1:0] n1579;
  wire [34-1:0] n158;
  wire [34-1:0] n1580;
  wire [34-1:0] n1581;
  wire [34-1:0] n1582;
  wire [34-1:0] n1583;
  wire [34-1:0] n1584;
  wire [34-1:0] n1585;
  wire [34-1:0] n1586;
  wire [34-1:0] n1587;
  wire [34-1:0] n1588;
  wire [34-1:0] n1589;
  wire [34-1:0] n159;
  wire [34-1:0] n1590;
  wire [34-1:0] n1591;
  wire [34-1:0] n1592;
  wire [34-1:0] n1593;
  wire [34-1:0] n1594;
  wire [34-1:0] n1595;
  wire [34-1:0] n1596;
  wire [34-1:0] n1597;
  wire [34-1:0] n1598;
  wire [34-1:0] n1599;
  wire [34-1:0] n16;
  wire [34-1:0] n160;
  wire [34-1:0] n1600;
  wire [34-1:0] n1601;
  wire [34-1:0] n1602;
  wire [34-1:0] n1603;
  wire [34-1:0] n1604;
  wire [34-1:0] n1605;
  wire [34-1:0] n1606;
  wire [34-1:0] n1607;
  wire [34-1:0] n1608;
  wire [34-1:0] n1609;
  wire [34-1:0] n161;
  wire [34-1:0] n1610;
  wire [34-1:0] n1611;
  wire [34-1:0] n1612;
  wire [34-1:0] n1613;
  wire [34-1:0] n1614;
  wire [34-1:0] n1615;
  wire [34-1:0] n1616;
  wire [34-1:0] n1617;
  wire [34-1:0] n1618;
  wire [34-1:0] n1619;
  wire [34-1:0] n162;
  wire [34-1:0] n1620;
  wire [34-1:0] n1621;
  wire [34-1:0] n1622;
  wire [34-1:0] n1623;
  wire [34-1:0] n1624;
  wire [34-1:0] n1625;
  wire [34-1:0] n1626;
  wire [34-1:0] n1627;
  wire [34-1:0] n1628;
  wire [34-1:0] n1629;
  wire [34-1:0] n163;
  wire [34-1:0] n1630;
  wire [34-1:0] n1631;
  wire [34-1:0] n1632;
  wire [34-1:0] n1633;
  wire [34-1:0] n1634;
  wire [34-1:0] n1635;
  wire [34-1:0] n1636;
  wire [34-1:0] n1637;
  wire [34-1:0] n1638;
  wire [34-1:0] n1639;
  wire [34-1:0] n164;
  wire [34-1:0] n1640;
  wire [34-1:0] n1641;
  wire [34-1:0] n1642;
  wire [34-1:0] n1643;
  wire [34-1:0] n1644;
  wire [34-1:0] n1645;
  wire [34-1:0] n1646;
  wire [34-1:0] n1647;
  wire [34-1:0] n1648;
  wire [34-1:0] n1649;
  wire [34-1:0] n165;
  wire [34-1:0] n1650;
  wire [34-1:0] n1651;
  wire [34-1:0] n1652;
  wire [34-1:0] n1653;
  wire [34-1:0] n1654;
  wire [34-1:0] n1655;
  wire [34-1:0] n1656;
  wire [34-1:0] n1657;
  wire [34-1:0] n1658;
  wire [34-1:0] n1659;
  wire [34-1:0] n166;
  wire [34-1:0] n1660;
  wire [34-1:0] n1661;
  wire [34-1:0] n1662;
  wire [34-1:0] n1663;
  wire [34-1:0] n1664;
  wire [34-1:0] n1665;
  wire [34-1:0] n1666;
  wire [34-1:0] n1667;
  wire [34-1:0] n1668;
  wire [34-1:0] n1669;
  wire [34-1:0] n167;
  wire [34-1:0] n1670;
  wire [34-1:0] n1671;
  wire [34-1:0] n1672;
  wire [34-1:0] n1673;
  wire [34-1:0] n1674;
  wire [34-1:0] n1675;
  wire [34-1:0] n1676;
  wire [34-1:0] n1677;
  wire [34-1:0] n1678;
  wire [34-1:0] n1679;
  wire [34-1:0] n168;
  wire [34-1:0] n1680;
  wire [34-1:0] n1681;
  wire [34-1:0] n1682;
  wire [34-1:0] n1683;
  wire [34-1:0] n1684;
  wire [34-1:0] n1685;
  wire [34-1:0] n1686;
  wire [34-1:0] n1687;
  wire [34-1:0] n1688;
  wire [34-1:0] n1689;
  wire [34-1:0] n169;
  wire [34-1:0] n1690;
  wire [34-1:0] n1691;
  wire [34-1:0] n1692;
  wire [34-1:0] n1693;
  wire [34-1:0] n1694;
  wire [34-1:0] n1695;
  wire [34-1:0] n1696;
  wire [34-1:0] n1697;
  wire [34-1:0] n1698;
  wire [34-1:0] n1699;
  wire [34-1:0] n17;
  wire [34-1:0] n170;
  wire [34-1:0] n1700;
  wire [34-1:0] n1701;
  wire [34-1:0] n1702;
  wire [34-1:0] n1703;
  wire [34-1:0] n1704;
  wire [34-1:0] n1705;
  wire [34-1:0] n1706;
  wire [34-1:0] n1707;
  wire [34-1:0] n1708;
  wire [34-1:0] n1709;
  wire [34-1:0] n171;
  wire [34-1:0] n1710;
  wire [34-1:0] n1711;
  wire [34-1:0] n1712;
  wire [34-1:0] n1713;
  wire [34-1:0] n1714;
  wire [34-1:0] n1715;
  wire [34-1:0] n1716;
  wire [34-1:0] n1717;
  wire [34-1:0] n1718;
  wire [34-1:0] n1719;
  wire [34-1:0] n172;
  wire [34-1:0] n1720;
  wire [34-1:0] n1721;
  wire [34-1:0] n1722;
  wire [34-1:0] n1723;
  wire [34-1:0] n1724;
  wire [34-1:0] n1725;
  wire [34-1:0] n1726;
  wire [34-1:0] n1727;
  wire [34-1:0] n1728;
  wire [34-1:0] n1729;
  wire [34-1:0] n173;
  wire [34-1:0] n1730;
  wire [34-1:0] n1731;
  wire [34-1:0] n1732;
  wire [34-1:0] n1733;
  wire [34-1:0] n1734;
  wire [34-1:0] n1735;
  wire [34-1:0] n1736;
  wire [34-1:0] n1737;
  wire [34-1:0] n1738;
  wire [34-1:0] n1739;
  wire [34-1:0] n174;
  wire [34-1:0] n1740;
  wire [34-1:0] n1741;
  wire [34-1:0] n1742;
  wire [34-1:0] n1743;
  wire [34-1:0] n1744;
  wire [34-1:0] n1745;
  wire [34-1:0] n1746;
  wire [34-1:0] n1747;
  wire [34-1:0] n1748;
  wire [34-1:0] n1749;
  wire [34-1:0] n175;
  wire [34-1:0] n1750;
  wire [34-1:0] n1751;
  wire [34-1:0] n1752;
  wire [34-1:0] n1753;
  wire [34-1:0] n1754;
  wire [34-1:0] n1755;
  wire [34-1:0] n1756;
  wire [34-1:0] n1757;
  wire [34-1:0] n1758;
  wire [34-1:0] n1759;
  wire [34-1:0] n176;
  wire [34-1:0] n1760;
  wire [34-1:0] n1761;
  wire [34-1:0] n1762;
  wire [34-1:0] n1763;
  wire [34-1:0] n1764;
  wire [34-1:0] n1765;
  wire [34-1:0] n1766;
  wire [34-1:0] n1767;
  wire [34-1:0] n1768;
  wire [34-1:0] n1769;
  wire [34-1:0] n177;
  wire [34-1:0] n1770;
  wire [34-1:0] n1771;
  wire [34-1:0] n1772;
  wire [34-1:0] n1773;
  wire [34-1:0] n1774;
  wire [34-1:0] n1775;
  wire [34-1:0] n1776;
  wire [34-1:0] n1777;
  wire [34-1:0] n1778;
  wire [34-1:0] n1779;
  wire [34-1:0] n178;
  wire [34-1:0] n1780;
  wire [34-1:0] n1781;
  wire [34-1:0] n1782;
  wire [34-1:0] n1783;
  wire [34-1:0] n1784;
  wire [34-1:0] n1785;
  wire [34-1:0] n1786;
  wire [34-1:0] n1787;
  wire [34-1:0] n1788;
  wire [34-1:0] n1789;
  wire [34-1:0] n179;
  wire [34-1:0] n1790;
  wire [34-1:0] n1791;
  wire [34-1:0] n1792;
  wire [34-1:0] n1793;
  wire [34-1:0] n1794;
  wire [34-1:0] n1795;
  wire [34-1:0] n1796;
  wire [34-1:0] n1797;
  wire [34-1:0] n1798;
  wire [34-1:0] n1799;
  wire [34-1:0] n18;
  wire [34-1:0] n180;
  wire [34-1:0] n1800;
  wire [34-1:0] n1801;
  wire [34-1:0] n1802;
  wire [34-1:0] n1803;
  wire [34-1:0] n1804;
  wire [34-1:0] n1805;
  wire [34-1:0] n1806;
  wire [34-1:0] n1807;
  wire [34-1:0] n1808;
  wire [34-1:0] n1809;
  wire [34-1:0] n181;
  wire [34-1:0] n1810;
  wire [34-1:0] n1811;
  wire [34-1:0] n1812;
  wire [34-1:0] n1813;
  wire [34-1:0] n1814;
  wire [34-1:0] n1815;
  wire [34-1:0] n1816;
  wire [34-1:0] n1817;
  wire [34-1:0] n1818;
  wire [34-1:0] n1819;
  wire [34-1:0] n182;
  wire [34-1:0] n1820;
  wire [34-1:0] n1821;
  wire [34-1:0] n1822;
  wire [34-1:0] n1823;
  wire [34-1:0] n1824;
  wire [34-1:0] n1825;
  wire [34-1:0] n1826;
  wire [34-1:0] n1827;
  wire [34-1:0] n1828;
  wire [34-1:0] n1829;
  wire [34-1:0] n183;
  wire [34-1:0] n1830;
  wire [34-1:0] n1831;
  wire [34-1:0] n1832;
  wire [34-1:0] n1833;
  wire [34-1:0] n1834;
  wire [34-1:0] n1835;
  wire [34-1:0] n1836;
  wire [34-1:0] n1837;
  wire [34-1:0] n1838;
  wire [34-1:0] n1839;
  wire [34-1:0] n184;
  wire [34-1:0] n1840;
  wire [34-1:0] n1841;
  wire [34-1:0] n1842;
  wire [34-1:0] n1843;
  wire [34-1:0] n1844;
  wire [34-1:0] n1845;
  wire [34-1:0] n1846;
  wire [34-1:0] n1847;
  wire [34-1:0] n1848;
  wire [34-1:0] n1849;
  wire [34-1:0] n185;
  wire [34-1:0] n1850;
  wire [34-1:0] n1851;
  wire [34-1:0] n1852;
  wire [34-1:0] n1853;
  wire [34-1:0] n1854;
  wire [34-1:0] n1855;
  wire [34-1:0] n1856;
  wire [34-1:0] n1857;
  wire [34-1:0] n1858;
  wire [34-1:0] n1859;
  wire [34-1:0] n186;
  wire [34-1:0] n1860;
  wire [34-1:0] n1861;
  wire [34-1:0] n1862;
  wire [34-1:0] n1863;
  wire [34-1:0] n1864;
  wire [34-1:0] n1865;
  wire [34-1:0] n1866;
  wire [34-1:0] n1867;
  wire [34-1:0] n1868;
  wire [34-1:0] n1869;
  wire [34-1:0] n187;
  wire [34-1:0] n1870;
  wire [34-1:0] n1871;
  wire [34-1:0] n1872;
  wire [34-1:0] n1873;
  wire [34-1:0] n1874;
  wire [34-1:0] n1875;
  wire [34-1:0] n1876;
  wire [34-1:0] n1877;
  wire [34-1:0] n1878;
  wire [34-1:0] n1879;
  wire [34-1:0] n188;
  wire [34-1:0] n1880;
  wire [34-1:0] n1881;
  wire [34-1:0] n1882;
  wire [34-1:0] n1883;
  wire [34-1:0] n1884;
  wire [34-1:0] n1885;
  wire [34-1:0] n1886;
  wire [34-1:0] n1887;
  wire [34-1:0] n1888;
  wire [34-1:0] n1889;
  wire [34-1:0] n189;
  wire [34-1:0] n1890;
  wire [34-1:0] n1891;
  wire [34-1:0] n1892;
  wire [34-1:0] n1893;
  wire [34-1:0] n1894;
  wire [34-1:0] n1895;
  wire [34-1:0] n1896;
  wire [34-1:0] n1897;
  wire [34-1:0] n1898;
  wire [34-1:0] n1899;
  wire [34-1:0] n19;
  wire [34-1:0] n190;
  wire [34-1:0] n1900;
  wire [34-1:0] n1901;
  wire [34-1:0] n1902;
  wire [34-1:0] n1903;
  wire [34-1:0] n1904;
  wire [34-1:0] n1905;
  wire [34-1:0] n1906;
  wire [34-1:0] n1907;
  wire [34-1:0] n1908;
  wire [34-1:0] n1909;
  wire [34-1:0] n191;
  wire [34-1:0] n1910;
  wire [34-1:0] n1911;
  wire [34-1:0] n1912;
  wire [34-1:0] n1913;
  wire [34-1:0] n1914;
  wire [34-1:0] n1915;
  wire [34-1:0] n1916;
  wire [34-1:0] n1917;
  wire [34-1:0] n1918;
  wire [34-1:0] n1919;
  wire [34-1:0] n192;
  wire [34-1:0] n1920;
  wire [34-1:0] n1921;
  wire [34-1:0] n1922;
  wire [34-1:0] n1923;
  wire [34-1:0] n1924;
  wire [34-1:0] n1925;
  wire [34-1:0] n1926;
  wire [34-1:0] n1927;
  wire [34-1:0] n1928;
  wire [34-1:0] n1929;
  wire [34-1:0] n193;
  wire [34-1:0] n1930;
  wire [34-1:0] n1931;
  wire [34-1:0] n1932;
  wire [34-1:0] n1933;
  wire [34-1:0] n1934;
  wire [34-1:0] n1935;
  wire [34-1:0] n1936;
  wire [34-1:0] n1937;
  wire [34-1:0] n1938;
  wire [34-1:0] n1939;
  wire [34-1:0] n194;
  wire [34-1:0] n1940;
  wire [34-1:0] n1941;
  wire [34-1:0] n1942;
  wire [34-1:0] n1943;
  wire [34-1:0] n1944;
  wire [34-1:0] n1945;
  wire [34-1:0] n1946;
  wire [34-1:0] n1947;
  wire [34-1:0] n1948;
  wire [34-1:0] n1949;
  wire [34-1:0] n195;
  wire [34-1:0] n1950;
  wire [34-1:0] n1951;
  wire [34-1:0] n1952;
  wire [34-1:0] n1953;
  wire [34-1:0] n1954;
  wire [34-1:0] n1955;
  wire [34-1:0] n1956;
  wire [34-1:0] n1957;
  wire [34-1:0] n1958;
  wire [34-1:0] n1959;
  wire [34-1:0] n196;
  wire [34-1:0] n1960;
  wire [34-1:0] n1961;
  wire [34-1:0] n1962;
  wire [34-1:0] n1963;
  wire [34-1:0] n1964;
  wire [34-1:0] n1965;
  wire [34-1:0] n1966;
  wire [34-1:0] n1967;
  wire [34-1:0] n1968;
  wire [34-1:0] n1969;
  wire [34-1:0] n197;
  wire [34-1:0] n1970;
  wire [34-1:0] n1971;
  wire [34-1:0] n1972;
  wire [34-1:0] n1973;
  wire [34-1:0] n1974;
  wire [34-1:0] n1975;
  wire [34-1:0] n1976;
  wire [34-1:0] n1977;
  wire [34-1:0] n1978;
  wire [34-1:0] n1979;
  wire [34-1:0] n198;
  wire [34-1:0] n1980;
  wire [34-1:0] n1981;
  wire [34-1:0] n1982;
  wire [34-1:0] n1983;
  wire [34-1:0] n1984;
  wire [34-1:0] n1985;
  wire [34-1:0] n1986;
  wire [34-1:0] n1987;
  wire [34-1:0] n1988;
  wire [34-1:0] n1989;
  wire [34-1:0] n199;
  wire [34-1:0] n1990;
  wire [34-1:0] n1991;
  wire [34-1:0] n1992;
  wire [34-1:0] n1993;
  wire [34-1:0] n1994;
  wire [34-1:0] n1995;
  wire [34-1:0] n1996;
  wire [34-1:0] n1997;
  wire [34-1:0] n1998;
  wire [34-1:0] n1999;
  wire [34-1:0] n2;
  wire [34-1:0] n20;
  wire [34-1:0] n200;
  wire [34-1:0] n2000;
  wire [34-1:0] n2001;
  wire [34-1:0] n2002;
  wire [34-1:0] n2003;
  wire [34-1:0] n2004;
  wire [34-1:0] n2005;
  wire [34-1:0] n2006;
  wire [34-1:0] n2007;
  wire [34-1:0] n2008;
  wire [34-1:0] n2009;
  wire [34-1:0] n201;
  wire [34-1:0] n2010;
  wire [34-1:0] n2011;
  wire [34-1:0] n2012;
  wire [34-1:0] n2013;
  wire [34-1:0] n2014;
  wire [34-1:0] n2015;
  wire [34-1:0] n2016;
  wire [34-1:0] n2017;
  wire [34-1:0] n2018;
  wire [34-1:0] n2019;
  wire [34-1:0] n202;
  wire [34-1:0] n2020;
  wire [34-1:0] n2021;
  wire [34-1:0] n2022;
  wire [34-1:0] n2023;
  wire [34-1:0] n2024;
  wire [34-1:0] n2025;
  wire [34-1:0] n2026;
  wire [34-1:0] n2027;
  wire [34-1:0] n2028;
  wire [34-1:0] n2029;
  wire [34-1:0] n203;
  wire [34-1:0] n2030;
  wire [34-1:0] n2031;
  wire [34-1:0] n2032;
  wire [34-1:0] n2033;
  wire [34-1:0] n2034;
  wire [34-1:0] n2035;
  wire [34-1:0] n2036;
  wire [34-1:0] n2037;
  wire [34-1:0] n2038;
  wire [34-1:0] n2039;
  wire [34-1:0] n204;
  wire [34-1:0] n2040;
  wire [34-1:0] n2041;
  wire [34-1:0] n2042;
  wire [34-1:0] n2043;
  wire [34-1:0] n2044;
  wire [34-1:0] n2045;
  wire [34-1:0] n2046;
  wire [34-1:0] n2047;
  wire [34-1:0] n2048;
  wire [34-1:0] n2049;
  wire [34-1:0] n205;
  wire [34-1:0] n2050;
  wire [34-1:0] n2051;
  wire [34-1:0] n2052;
  wire [34-1:0] n2053;
  wire [34-1:0] n2054;
  wire [34-1:0] n2055;
  wire [34-1:0] n2056;
  wire [34-1:0] n2057;
  wire [34-1:0] n2058;
  wire [34-1:0] n2059;
  wire [34-1:0] n206;
  wire [34-1:0] n2060;
  wire [34-1:0] n2061;
  wire [34-1:0] n2062;
  wire [34-1:0] n2063;
  wire [34-1:0] n2064;
  wire [34-1:0] n2065;
  wire [34-1:0] n2066;
  wire [34-1:0] n2067;
  wire [34-1:0] n2068;
  wire [34-1:0] n2069;
  wire [34-1:0] n207;
  wire [34-1:0] n2070;
  wire [34-1:0] n2071;
  wire [34-1:0] n2072;
  wire [34-1:0] n2073;
  wire [34-1:0] n2074;
  wire [34-1:0] n2075;
  wire [34-1:0] n2076;
  wire [34-1:0] n2077;
  wire [34-1:0] n2078;
  wire [34-1:0] n2079;
  wire [34-1:0] n208;
  wire [34-1:0] n2080;
  wire [34-1:0] n2081;
  wire [34-1:0] n2082;
  wire [34-1:0] n2083;
  wire [34-1:0] n2084;
  wire [34-1:0] n2085;
  wire [34-1:0] n2086;
  wire [34-1:0] n2087;
  wire [34-1:0] n2088;
  wire [34-1:0] n2089;
  wire [34-1:0] n209;
  wire [34-1:0] n2090;
  wire [34-1:0] n2091;
  wire [34-1:0] n2092;
  wire [34-1:0] n2093;
  wire [34-1:0] n2094;
  wire [34-1:0] n2095;
  wire [34-1:0] n2096;
  wire [34-1:0] n2097;
  wire [34-1:0] n2098;
  wire [34-1:0] n2099;
  wire [34-1:0] n21;
  wire [34-1:0] n210;
  wire [34-1:0] n2100;
  wire [34-1:0] n2101;
  wire [34-1:0] n2102;
  wire [34-1:0] n2103;
  wire [34-1:0] n2104;
  wire [34-1:0] n2105;
  wire [34-1:0] n2106;
  wire [34-1:0] n2107;
  wire [34-1:0] n2108;
  wire [34-1:0] n2109;
  wire [34-1:0] n211;
  wire [34-1:0] n2110;
  wire [34-1:0] n2111;
  wire [34-1:0] n2112;
  wire [34-1:0] n2113;
  wire [34-1:0] n2114;
  wire [34-1:0] n2115;
  wire [34-1:0] n2116;
  wire [34-1:0] n2117;
  wire [34-1:0] n2118;
  wire [34-1:0] n2119;
  wire [34-1:0] n212;
  wire [34-1:0] n2120;
  wire [34-1:0] n2121;
  wire [34-1:0] n2122;
  wire [34-1:0] n2123;
  wire [34-1:0] n2124;
  wire [34-1:0] n2125;
  wire [34-1:0] n2126;
  wire [34-1:0] n2127;
  wire [34-1:0] n2128;
  wire [34-1:0] n2129;
  wire [34-1:0] n213;
  wire [34-1:0] n2130;
  wire [34-1:0] n2131;
  wire [34-1:0] n2132;
  wire [34-1:0] n2133;
  wire [34-1:0] n2134;
  wire [34-1:0] n2135;
  wire [34-1:0] n2136;
  wire [34-1:0] n2137;
  wire [34-1:0] n2138;
  wire [34-1:0] n2139;
  wire [34-1:0] n214;
  wire [34-1:0] n2140;
  wire [34-1:0] n2141;
  wire [34-1:0] n2142;
  wire [34-1:0] n2143;
  wire [34-1:0] n2144;
  wire [34-1:0] n2145;
  wire [34-1:0] n2146;
  wire [34-1:0] n2147;
  wire [34-1:0] n2148;
  wire [34-1:0] n2149;
  wire [34-1:0] n215;
  wire [34-1:0] n2150;
  wire [34-1:0] n2151;
  wire [34-1:0] n2152;
  wire [34-1:0] n2153;
  wire [34-1:0] n2154;
  wire [34-1:0] n2155;
  wire [34-1:0] n2156;
  wire [34-1:0] n2157;
  wire [34-1:0] n2158;
  wire [34-1:0] n2159;
  wire [34-1:0] n216;
  wire [34-1:0] n2160;
  wire [34-1:0] n2161;
  wire [34-1:0] n2162;
  wire [34-1:0] n2163;
  wire [34-1:0] n2164;
  wire [34-1:0] n2165;
  wire [34-1:0] n2166;
  wire [34-1:0] n2167;
  wire [34-1:0] n2168;
  wire [34-1:0] n2169;
  wire [34-1:0] n217;
  wire [34-1:0] n2170;
  wire [34-1:0] n2171;
  wire [34-1:0] n2172;
  wire [34-1:0] n2173;
  wire [34-1:0] n2174;
  wire [34-1:0] n2175;
  wire [34-1:0] n2176;
  wire [34-1:0] n2177;
  wire [34-1:0] n2178;
  wire [34-1:0] n2179;
  wire [34-1:0] n218;
  wire [34-1:0] n2180;
  wire [34-1:0] n2181;
  wire [34-1:0] n2182;
  wire [34-1:0] n2183;
  wire [34-1:0] n2184;
  wire [34-1:0] n2185;
  wire [34-1:0] n2186;
  wire [34-1:0] n2187;
  wire [34-1:0] n2188;
  wire [34-1:0] n2189;
  wire [34-1:0] n219;
  wire [34-1:0] n2190;
  wire [34-1:0] n2191;
  wire [34-1:0] n2192;
  wire [34-1:0] n2193;
  wire [34-1:0] n2194;
  wire [34-1:0] n2195;
  wire [34-1:0] n2196;
  wire [34-1:0] n2197;
  wire [34-1:0] n2198;
  wire [34-1:0] n2199;
  wire [34-1:0] n22;
  wire [34-1:0] n220;
  wire [34-1:0] n2200;
  wire [34-1:0] n2201;
  wire [34-1:0] n2202;
  wire [34-1:0] n2203;
  wire [34-1:0] n2204;
  wire [34-1:0] n2205;
  wire [34-1:0] n2206;
  wire [34-1:0] n2207;
  wire [34-1:0] n2208;
  wire [34-1:0] n2209;
  wire [34-1:0] n221;
  wire [34-1:0] n2210;
  wire [34-1:0] n2211;
  wire [34-1:0] n2212;
  wire [34-1:0] n2213;
  wire [34-1:0] n2214;
  wire [34-1:0] n2215;
  wire [34-1:0] n2216;
  wire [34-1:0] n2217;
  wire [34-1:0] n2218;
  wire [34-1:0] n2219;
  wire [34-1:0] n222;
  wire [34-1:0] n2220;
  wire [34-1:0] n2221;
  wire [34-1:0] n2222;
  wire [34-1:0] n2223;
  wire [34-1:0] n2224;
  wire [34-1:0] n2225;
  wire [34-1:0] n2226;
  wire [34-1:0] n2227;
  wire [34-1:0] n2228;
  wire [34-1:0] n2229;
  wire [34-1:0] n223;
  wire [34-1:0] n2230;
  wire [34-1:0] n2231;
  wire [34-1:0] n2232;
  wire [34-1:0] n2233;
  wire [34-1:0] n2234;
  wire [34-1:0] n2235;
  wire [34-1:0] n2236;
  wire [34-1:0] n2237;
  wire [34-1:0] n2238;
  wire [34-1:0] n2239;
  wire [34-1:0] n224;
  wire [34-1:0] n2240;
  wire [34-1:0] n2241;
  wire [34-1:0] n2242;
  wire [34-1:0] n2243;
  wire [34-1:0] n2244;
  wire [34-1:0] n2245;
  wire [34-1:0] n2246;
  wire [34-1:0] n2247;
  wire [34-1:0] n2248;
  wire [34-1:0] n2249;
  wire [34-1:0] n225;
  wire [34-1:0] n2250;
  wire [34-1:0] n2251;
  wire [34-1:0] n2252;
  wire [34-1:0] n2253;
  wire [34-1:0] n2254;
  wire [34-1:0] n2255;
  wire [34-1:0] n2256;
  wire [34-1:0] n2257;
  wire [34-1:0] n2258;
  wire [34-1:0] n2259;
  wire [34-1:0] n226;
  wire [34-1:0] n2260;
  wire [34-1:0] n2261;
  wire [34-1:0] n2262;
  wire [34-1:0] n2263;
  wire [34-1:0] n2264;
  wire [34-1:0] n2265;
  wire [34-1:0] n2266;
  wire [34-1:0] n2267;
  wire [34-1:0] n2268;
  wire [34-1:0] n2269;
  wire [34-1:0] n227;
  wire [34-1:0] n2270;
  wire [34-1:0] n2271;
  wire [34-1:0] n2272;
  wire [34-1:0] n2273;
  wire [34-1:0] n2274;
  wire [34-1:0] n2275;
  wire [34-1:0] n2276;
  wire [34-1:0] n2277;
  wire [34-1:0] n2278;
  wire [34-1:0] n2279;
  wire [34-1:0] n228;
  wire [34-1:0] n2280;
  wire [34-1:0] n2281;
  wire [34-1:0] n2282;
  wire [34-1:0] n2283;
  wire [34-1:0] n2284;
  wire [34-1:0] n2285;
  wire [34-1:0] n2286;
  wire [34-1:0] n2287;
  wire [34-1:0] n2288;
  wire [34-1:0] n2289;
  wire [34-1:0] n229;
  wire [34-1:0] n2290;
  wire [34-1:0] n2291;
  wire [34-1:0] n2292;
  wire [34-1:0] n2293;
  wire [34-1:0] n2294;
  wire [34-1:0] n2295;
  wire [34-1:0] n2296;
  wire [34-1:0] n2297;
  wire [34-1:0] n2298;
  wire [34-1:0] n2299;
  wire [34-1:0] n23;
  wire [34-1:0] n230;
  wire [34-1:0] n2300;
  wire [34-1:0] n2301;
  wire [34-1:0] n2302;
  wire [34-1:0] n2303;
  wire [34-1:0] n2304;
  wire [34-1:0] n2305;
  wire [34-1:0] n2306;
  wire [34-1:0] n2307;
  wire [34-1:0] n2308;
  wire [34-1:0] n2309;
  wire [34-1:0] n231;
  wire [34-1:0] n2310;
  wire [34-1:0] n2311;
  wire [34-1:0] n2312;
  wire [34-1:0] n2313;
  wire [34-1:0] n2314;
  wire [34-1:0] n2315;
  wire [34-1:0] n2316;
  wire [34-1:0] n2317;
  wire [34-1:0] n2318;
  wire [34-1:0] n2319;
  wire [34-1:0] n232;
  wire [34-1:0] n2320;
  wire [34-1:0] n2321;
  wire [34-1:0] n2322;
  wire [34-1:0] n2323;
  wire [34-1:0] n2324;
  wire [34-1:0] n2325;
  wire [34-1:0] n2326;
  wire [34-1:0] n2327;
  wire [34-1:0] n2328;
  wire [34-1:0] n2329;
  wire [34-1:0] n233;
  wire [34-1:0] n2330;
  wire [34-1:0] n2331;
  wire [34-1:0] n2332;
  wire [34-1:0] n2333;
  wire [34-1:0] n2334;
  wire [34-1:0] n2335;
  wire [34-1:0] n2336;
  wire [34-1:0] n2337;
  wire [34-1:0] n2338;
  wire [34-1:0] n2339;
  wire [34-1:0] n234;
  wire [34-1:0] n2340;
  wire [34-1:0] n2341;
  wire [34-1:0] n2342;
  wire [34-1:0] n2343;
  wire [34-1:0] n2344;
  wire [34-1:0] n2345;
  wire [34-1:0] n2346;
  wire [34-1:0] n2347;
  wire [34-1:0] n2348;
  wire [34-1:0] n2349;
  wire [34-1:0] n235;
  wire [34-1:0] n2350;
  wire [34-1:0] n2351;
  wire [34-1:0] n2352;
  wire [34-1:0] n2353;
  wire [34-1:0] n2354;
  wire [34-1:0] n2355;
  wire [34-1:0] n2356;
  wire [34-1:0] n2357;
  wire [34-1:0] n2358;
  wire [34-1:0] n2359;
  wire [34-1:0] n236;
  wire [34-1:0] n2360;
  wire [34-1:0] n2361;
  wire [34-1:0] n2362;
  wire [34-1:0] n2363;
  wire [34-1:0] n2364;
  wire [34-1:0] n2365;
  wire [34-1:0] n2366;
  wire [34-1:0] n2367;
  wire [34-1:0] n2368;
  wire [34-1:0] n2369;
  wire [34-1:0] n237;
  wire [34-1:0] n2370;
  wire [34-1:0] n2371;
  wire [34-1:0] n2372;
  wire [34-1:0] n2373;
  wire [34-1:0] n2374;
  wire [34-1:0] n2375;
  wire [34-1:0] n2376;
  wire [34-1:0] n2377;
  wire [34-1:0] n2378;
  wire [34-1:0] n2379;
  wire [34-1:0] n238;
  wire [34-1:0] n2380;
  wire [34-1:0] n2381;
  wire [34-1:0] n2382;
  wire [34-1:0] n2383;
  wire [34-1:0] n2384;
  wire [34-1:0] n2385;
  wire [34-1:0] n2386;
  wire [34-1:0] n2387;
  wire [34-1:0] n2388;
  wire [34-1:0] n2389;
  wire [34-1:0] n239;
  wire [34-1:0] n2390;
  wire [34-1:0] n2391;
  wire [34-1:0] n2392;
  wire [34-1:0] n2393;
  wire [34-1:0] n2394;
  wire [34-1:0] n2395;
  wire [34-1:0] n2396;
  wire [34-1:0] n2397;
  wire [34-1:0] n2398;
  wire [34-1:0] n2399;
  wire [34-1:0] n24;
  wire [34-1:0] n240;
  wire [34-1:0] n2400;
  wire [34-1:0] n2401;
  wire [34-1:0] n2402;
  wire [34-1:0] n2403;
  wire [34-1:0] n2404;
  wire [34-1:0] n2405;
  wire [34-1:0] n2406;
  wire [34-1:0] n2407;
  wire [34-1:0] n2408;
  wire [34-1:0] n2409;
  wire [34-1:0] n241;
  wire [34-1:0] n2410;
  wire [34-1:0] n2411;
  wire [34-1:0] n2412;
  wire [34-1:0] n2413;
  wire [34-1:0] n2414;
  wire [34-1:0] n2415;
  wire [34-1:0] n2416;
  wire [34-1:0] n2417;
  wire [34-1:0] n2418;
  wire [34-1:0] n2419;
  wire [34-1:0] n242;
  wire [34-1:0] n2420;
  wire [34-1:0] n2421;
  wire [34-1:0] n2422;
  wire [34-1:0] n2423;
  wire [34-1:0] n2424;
  wire [34-1:0] n2425;
  wire [34-1:0] n2426;
  wire [34-1:0] n2427;
  wire [34-1:0] n2428;
  wire [34-1:0] n2429;
  wire [34-1:0] n243;
  wire [34-1:0] n2430;
  wire [34-1:0] n2431;
  wire [34-1:0] n2432;
  wire [34-1:0] n2433;
  wire [34-1:0] n2434;
  wire [34-1:0] n2435;
  wire [34-1:0] n2436;
  wire [34-1:0] n2437;
  wire [34-1:0] n2438;
  wire [34-1:0] n2439;
  wire [34-1:0] n244;
  wire [34-1:0] n2440;
  wire [34-1:0] n2441;
  wire [34-1:0] n2442;
  wire [34-1:0] n2443;
  wire [34-1:0] n2444;
  wire [34-1:0] n2445;
  wire [34-1:0] n2446;
  wire [34-1:0] n2447;
  wire [34-1:0] n2448;
  wire [34-1:0] n2449;
  wire [34-1:0] n245;
  wire [34-1:0] n246;
  wire [34-1:0] n247;
  wire [34-1:0] n248;
  wire [34-1:0] n249;
  wire [34-1:0] n25;
  wire [34-1:0] n250;
  wire [34-1:0] n251;
  wire [34-1:0] n252;
  wire [34-1:0] n253;
  wire [34-1:0] n254;
  wire [34-1:0] n255;
  wire [34-1:0] n256;
  wire [34-1:0] n257;
  wire [34-1:0] n258;
  wire [34-1:0] n259;
  wire [34-1:0] n26;
  wire [34-1:0] n260;
  wire [34-1:0] n261;
  wire [34-1:0] n262;
  wire [34-1:0] n263;
  wire [34-1:0] n264;
  wire [34-1:0] n265;
  wire [34-1:0] n266;
  wire [34-1:0] n267;
  wire [34-1:0] n268;
  wire [34-1:0] n269;
  wire [34-1:0] n27;
  wire [34-1:0] n270;
  wire [34-1:0] n271;
  wire [34-1:0] n272;
  wire [34-1:0] n273;
  wire [34-1:0] n274;
  wire [34-1:0] n275;
  wire [34-1:0] n276;
  wire [34-1:0] n277;
  wire [34-1:0] n278;
  wire [34-1:0] n279;
  wire [34-1:0] n28;
  wire [34-1:0] n280;
  wire [34-1:0] n281;
  wire [34-1:0] n282;
  wire [34-1:0] n283;
  wire [34-1:0] n284;
  wire [34-1:0] n285;
  wire [34-1:0] n286;
  wire [34-1:0] n287;
  wire [34-1:0] n288;
  wire [34-1:0] n289;
  wire [34-1:0] n29;
  wire [34-1:0] n290;
  wire [34-1:0] n291;
  wire [34-1:0] n292;
  wire [34-1:0] n293;
  wire [34-1:0] n294;
  wire [34-1:0] n295;
  wire [34-1:0] n296;
  wire [34-1:0] n297;
  wire [34-1:0] n298;
  wire [34-1:0] n299;
  wire [34-1:0] n3;
  wire [34-1:0] n30;
  wire [34-1:0] n300;
  wire [34-1:0] n301;
  wire [34-1:0] n302;
  wire [34-1:0] n303;
  wire [34-1:0] n304;
  wire [34-1:0] n305;
  wire [34-1:0] n306;
  wire [34-1:0] n307;
  wire [34-1:0] n308;
  wire [34-1:0] n309;
  wire [34-1:0] n31;
  wire [34-1:0] n310;
  wire [34-1:0] n311;
  wire [34-1:0] n312;
  wire [34-1:0] n313;
  wire [34-1:0] n314;
  wire [34-1:0] n315;
  wire [34-1:0] n316;
  wire [34-1:0] n317;
  wire [34-1:0] n318;
  wire [34-1:0] n319;
  wire [34-1:0] n32;
  wire [34-1:0] n320;
  wire [34-1:0] n321;
  wire [34-1:0] n322;
  wire [34-1:0] n323;
  wire [34-1:0] n324;
  wire [34-1:0] n325;
  wire [34-1:0] n326;
  wire [34-1:0] n327;
  wire [34-1:0] n328;
  wire [34-1:0] n329;
  wire [34-1:0] n33;
  wire [34-1:0] n330;
  wire [34-1:0] n331;
  wire [34-1:0] n332;
  wire [34-1:0] n333;
  wire [34-1:0] n334;
  wire [34-1:0] n335;
  wire [34-1:0] n336;
  wire [34-1:0] n337;
  wire [34-1:0] n338;
  wire [34-1:0] n339;
  wire [34-1:0] n34;
  wire [34-1:0] n340;
  wire [34-1:0] n341;
  wire [34-1:0] n342;
  wire [34-1:0] n343;
  wire [34-1:0] n344;
  wire [34-1:0] n345;
  wire [34-1:0] n346;
  wire [34-1:0] n347;
  wire [34-1:0] n348;
  wire [34-1:0] n349;
  wire [34-1:0] n35;
  wire [34-1:0] n350;
  wire [34-1:0] n351;
  wire [34-1:0] n352;
  wire [34-1:0] n353;
  wire [34-1:0] n354;
  wire [34-1:0] n355;
  wire [34-1:0] n356;
  wire [34-1:0] n357;
  wire [34-1:0] n358;
  wire [34-1:0] n359;
  wire [34-1:0] n36;
  wire [34-1:0] n360;
  wire [34-1:0] n361;
  wire [34-1:0] n362;
  wire [34-1:0] n363;
  wire [34-1:0] n364;
  wire [34-1:0] n365;
  wire [34-1:0] n366;
  wire [34-1:0] n367;
  wire [34-1:0] n368;
  wire [34-1:0] n369;
  wire [34-1:0] n37;
  wire [34-1:0] n370;
  wire [34-1:0] n371;
  wire [34-1:0] n372;
  wire [34-1:0] n373;
  wire [34-1:0] n374;
  wire [34-1:0] n375;
  wire [34-1:0] n376;
  wire [34-1:0] n377;
  wire [34-1:0] n378;
  wire [34-1:0] n379;
  wire [34-1:0] n38;
  wire [34-1:0] n380;
  wire [34-1:0] n381;
  wire [34-1:0] n382;
  wire [34-1:0] n383;
  wire [34-1:0] n384;
  wire [34-1:0] n385;
  wire [34-1:0] n386;
  wire [34-1:0] n387;
  wire [34-1:0] n388;
  wire [34-1:0] n389;
  wire [34-1:0] n39;
  wire [34-1:0] n390;
  wire [34-1:0] n391;
  wire [34-1:0] n392;
  wire [34-1:0] n393;
  wire [34-1:0] n394;
  wire [34-1:0] n395;
  wire [34-1:0] n396;
  wire [34-1:0] n397;
  wire [34-1:0] n398;
  wire [34-1:0] n399;
  wire [34-1:0] n4;
  wire [34-1:0] n40;
  wire [34-1:0] n400;
  wire [34-1:0] n401;
  wire [34-1:0] n402;
  wire [34-1:0] n403;
  wire [34-1:0] n404;
  wire [34-1:0] n405;
  wire [34-1:0] n406;
  wire [34-1:0] n407;
  wire [34-1:0] n408;
  wire [34-1:0] n409;
  wire [34-1:0] n41;
  wire [34-1:0] n410;
  wire [34-1:0] n411;
  wire [34-1:0] n412;
  wire [34-1:0] n413;
  wire [34-1:0] n414;
  wire [34-1:0] n415;
  wire [34-1:0] n416;
  wire [34-1:0] n417;
  wire [34-1:0] n418;
  wire [34-1:0] n419;
  wire [34-1:0] n42;
  wire [34-1:0] n420;
  wire [34-1:0] n421;
  wire [34-1:0] n422;
  wire [34-1:0] n423;
  wire [34-1:0] n424;
  wire [34-1:0] n425;
  wire [34-1:0] n426;
  wire [34-1:0] n427;
  wire [34-1:0] n428;
  wire [34-1:0] n429;
  wire [34-1:0] n43;
  wire [34-1:0] n430;
  wire [34-1:0] n431;
  wire [34-1:0] n432;
  wire [34-1:0] n433;
  wire [34-1:0] n434;
  wire [34-1:0] n435;
  wire [34-1:0] n436;
  wire [34-1:0] n437;
  wire [34-1:0] n438;
  wire [34-1:0] n439;
  wire [34-1:0] n44;
  wire [34-1:0] n440;
  wire [34-1:0] n441;
  wire [34-1:0] n442;
  wire [34-1:0] n443;
  wire [34-1:0] n444;
  wire [34-1:0] n445;
  wire [34-1:0] n446;
  wire [34-1:0] n447;
  wire [34-1:0] n448;
  wire [34-1:0] n449;
  wire [34-1:0] n45;
  wire [34-1:0] n450;
  wire [34-1:0] n451;
  wire [34-1:0] n452;
  wire [34-1:0] n453;
  wire [34-1:0] n454;
  wire [34-1:0] n455;
  wire [34-1:0] n456;
  wire [34-1:0] n457;
  wire [34-1:0] n458;
  wire [34-1:0] n459;
  wire [34-1:0] n46;
  wire [34-1:0] n460;
  wire [34-1:0] n461;
  wire [34-1:0] n462;
  wire [34-1:0] n463;
  wire [34-1:0] n464;
  wire [34-1:0] n465;
  wire [34-1:0] n466;
  wire [34-1:0] n467;
  wire [34-1:0] n468;
  wire [34-1:0] n469;
  wire [34-1:0] n47;
  wire [34-1:0] n470;
  wire [34-1:0] n471;
  wire [34-1:0] n472;
  wire [34-1:0] n473;
  wire [34-1:0] n474;
  wire [34-1:0] n475;
  wire [34-1:0] n476;
  wire [34-1:0] n477;
  wire [34-1:0] n478;
  wire [34-1:0] n479;
  wire [34-1:0] n48;
  wire [34-1:0] n480;
  wire [34-1:0] n481;
  wire [34-1:0] n482;
  wire [34-1:0] n483;
  wire [34-1:0] n484;
  wire [34-1:0] n485;
  wire [34-1:0] n486;
  wire [34-1:0] n487;
  wire [34-1:0] n488;
  wire [34-1:0] n489;
  wire [34-1:0] n49;
  wire [34-1:0] n490;
  wire [34-1:0] n491;
  wire [34-1:0] n492;
  wire [34-1:0] n493;
  wire [34-1:0] n494;
  wire [34-1:0] n495;
  wire [34-1:0] n496;
  wire [34-1:0] n497;
  wire [34-1:0] n498;
  wire [34-1:0] n499;
  wire [34-1:0] n5;
  wire [34-1:0] n50;
  wire [34-1:0] n500;
  wire [34-1:0] n501;
  wire [34-1:0] n502;
  wire [34-1:0] n503;
  wire [34-1:0] n504;
  wire [34-1:0] n505;
  wire [34-1:0] n506;
  wire [34-1:0] n507;
  wire [34-1:0] n508;
  wire [34-1:0] n509;
  wire [34-1:0] n51;
  wire [34-1:0] n510;
  wire [34-1:0] n511;
  wire [34-1:0] n512;
  wire [34-1:0] n513;
  wire [34-1:0] n514;
  wire [34-1:0] n515;
  wire [34-1:0] n516;
  wire [34-1:0] n517;
  wire [34-1:0] n518;
  wire [34-1:0] n519;
  wire [34-1:0] n52;
  wire [34-1:0] n520;
  wire [34-1:0] n521;
  wire [34-1:0] n522;
  wire [34-1:0] n523;
  wire [34-1:0] n524;
  wire [34-1:0] n525;
  wire [34-1:0] n526;
  wire [34-1:0] n527;
  wire [34-1:0] n528;
  wire [34-1:0] n529;
  wire [34-1:0] n53;
  wire [34-1:0] n530;
  wire [34-1:0] n531;
  wire [34-1:0] n532;
  wire [34-1:0] n533;
  wire [34-1:0] n534;
  wire [34-1:0] n535;
  wire [34-1:0] n536;
  wire [34-1:0] n537;
  wire [34-1:0] n538;
  wire [34-1:0] n539;
  wire [34-1:0] n54;
  wire [34-1:0] n540;
  wire [34-1:0] n541;
  wire [34-1:0] n542;
  wire [34-1:0] n543;
  wire [34-1:0] n544;
  wire [34-1:0] n545;
  wire [34-1:0] n546;
  wire [34-1:0] n547;
  wire [34-1:0] n548;
  wire [34-1:0] n549;
  wire [34-1:0] n55;
  wire [34-1:0] n550;
  wire [34-1:0] n551;
  wire [34-1:0] n552;
  wire [34-1:0] n553;
  wire [34-1:0] n554;
  wire [34-1:0] n555;
  wire [34-1:0] n556;
  wire [34-1:0] n557;
  wire [34-1:0] n558;
  wire [34-1:0] n559;
  wire [34-1:0] n56;
  wire [34-1:0] n560;
  wire [34-1:0] n561;
  wire [34-1:0] n562;
  wire [34-1:0] n563;
  wire [34-1:0] n564;
  wire [34-1:0] n565;
  wire [34-1:0] n566;
  wire [34-1:0] n567;
  wire [34-1:0] n568;
  wire [34-1:0] n569;
  wire [34-1:0] n57;
  wire [34-1:0] n570;
  wire [34-1:0] n571;
  wire [34-1:0] n572;
  wire [34-1:0] n573;
  wire [34-1:0] n574;
  wire [34-1:0] n575;
  wire [34-1:0] n576;
  wire [34-1:0] n577;
  wire [34-1:0] n578;
  wire [34-1:0] n579;
  wire [34-1:0] n58;
  wire [34-1:0] n580;
  wire [34-1:0] n581;
  wire [34-1:0] n582;
  wire [34-1:0] n583;
  wire [34-1:0] n584;
  wire [34-1:0] n585;
  wire [34-1:0] n586;
  wire [34-1:0] n587;
  wire [34-1:0] n588;
  wire [34-1:0] n589;
  wire [34-1:0] n59;
  wire [34-1:0] n590;
  wire [34-1:0] n591;
  wire [34-1:0] n592;
  wire [34-1:0] n593;
  wire [34-1:0] n594;
  wire [34-1:0] n595;
  wire [34-1:0] n596;
  wire [34-1:0] n597;
  wire [34-1:0] n598;
  wire [34-1:0] n599;
  wire [34-1:0] n6;
  wire [34-1:0] n60;
  wire [34-1:0] n600;
  wire [34-1:0] n601;
  wire [34-1:0] n602;
  wire [34-1:0] n603;
  wire [34-1:0] n604;
  wire [34-1:0] n605;
  wire [34-1:0] n606;
  wire [34-1:0] n607;
  wire [34-1:0] n608;
  wire [34-1:0] n609;
  wire [34-1:0] n61;
  wire [34-1:0] n610;
  wire [34-1:0] n611;
  wire [34-1:0] n612;
  wire [34-1:0] n613;
  wire [34-1:0] n614;
  wire [34-1:0] n615;
  wire [34-1:0] n616;
  wire [34-1:0] n617;
  wire [34-1:0] n618;
  wire [34-1:0] n619;
  wire [34-1:0] n62;
  wire [34-1:0] n620;
  wire [34-1:0] n621;
  wire [34-1:0] n622;
  wire [34-1:0] n623;
  wire [34-1:0] n624;
  wire [34-1:0] n625;
  wire [34-1:0] n626;
  wire [34-1:0] n627;
  wire [34-1:0] n628;
  wire [34-1:0] n629;
  wire [34-1:0] n63;
  wire [34-1:0] n630;
  wire [34-1:0] n631;
  wire [34-1:0] n632;
  wire [34-1:0] n633;
  wire [34-1:0] n634;
  wire [34-1:0] n635;
  wire [34-1:0] n636;
  wire [34-1:0] n637;
  wire [34-1:0] n638;
  wire [34-1:0] n639;
  wire [34-1:0] n64;
  wire [34-1:0] n640;
  wire [34-1:0] n641;
  wire [34-1:0] n642;
  wire [34-1:0] n643;
  wire [34-1:0] n644;
  wire [34-1:0] n645;
  wire [34-1:0] n646;
  wire [34-1:0] n647;
  wire [34-1:0] n648;
  wire [34-1:0] n649;
  wire [34-1:0] n65;
  wire [34-1:0] n650;
  wire [34-1:0] n651;
  wire [34-1:0] n652;
  wire [34-1:0] n653;
  wire [34-1:0] n654;
  wire [34-1:0] n655;
  wire [34-1:0] n656;
  wire [34-1:0] n657;
  wire [34-1:0] n658;
  wire [34-1:0] n659;
  wire [34-1:0] n66;
  wire [34-1:0] n660;
  wire [34-1:0] n661;
  wire [34-1:0] n662;
  wire [34-1:0] n663;
  wire [34-1:0] n664;
  wire [34-1:0] n665;
  wire [34-1:0] n666;
  wire [34-1:0] n667;
  wire [34-1:0] n668;
  wire [34-1:0] n669;
  wire [34-1:0] n67;
  wire [34-1:0] n670;
  wire [34-1:0] n671;
  wire [34-1:0] n672;
  wire [34-1:0] n673;
  wire [34-1:0] n674;
  wire [34-1:0] n675;
  wire [34-1:0] n676;
  wire [34-1:0] n677;
  wire [34-1:0] n678;
  wire [34-1:0] n679;
  wire [34-1:0] n68;
  wire [34-1:0] n680;
  wire [34-1:0] n681;
  wire [34-1:0] n682;
  wire [34-1:0] n683;
  wire [34-1:0] n684;
  wire [34-1:0] n685;
  wire [34-1:0] n686;
  wire [34-1:0] n687;
  wire [34-1:0] n688;
  wire [34-1:0] n689;
  wire [34-1:0] n69;
  wire [34-1:0] n690;
  wire [34-1:0] n691;
  wire [34-1:0] n692;
  wire [34-1:0] n693;
  wire [34-1:0] n694;
  wire [34-1:0] n695;
  wire [34-1:0] n696;
  wire [34-1:0] n697;
  wire [34-1:0] n698;
  wire [34-1:0] n699;
  wire [34-1:0] n7;
  wire [34-1:0] n70;
  wire [34-1:0] n700;
  wire [34-1:0] n701;
  wire [34-1:0] n702;
  wire [34-1:0] n703;
  wire [34-1:0] n704;
  wire [34-1:0] n705;
  wire [34-1:0] n706;
  wire [34-1:0] n707;
  wire [34-1:0] n708;
  wire [34-1:0] n709;
  wire [34-1:0] n71;
  wire [34-1:0] n710;
  wire [34-1:0] n711;
  wire [34-1:0] n712;
  wire [34-1:0] n713;
  wire [34-1:0] n714;
  wire [34-1:0] n715;
  wire [34-1:0] n716;
  wire [34-1:0] n717;
  wire [34-1:0] n718;
  wire [34-1:0] n719;
  wire [34-1:0] n72;
  wire [34-1:0] n720;
  wire [34-1:0] n721;
  wire [34-1:0] n722;
  wire [34-1:0] n723;
  wire [34-1:0] n724;
  wire [34-1:0] n725;
  wire [34-1:0] n726;
  wire [34-1:0] n727;
  wire [34-1:0] n728;
  wire [34-1:0] n729;
  wire [34-1:0] n73;
  wire [34-1:0] n730;
  wire [34-1:0] n731;
  wire [34-1:0] n732;
  wire [34-1:0] n733;
  wire [34-1:0] n734;
  wire [34-1:0] n735;
  wire [34-1:0] n736;
  wire [34-1:0] n737;
  wire [34-1:0] n738;
  wire [34-1:0] n739;
  wire [34-1:0] n74;
  wire [34-1:0] n740;
  wire [34-1:0] n741;
  wire [34-1:0] n742;
  wire [34-1:0] n743;
  wire [34-1:0] n744;
  wire [34-1:0] n745;
  wire [34-1:0] n746;
  wire [34-1:0] n747;
  wire [34-1:0] n748;
  wire [34-1:0] n749;
  wire [34-1:0] n75;
  wire [34-1:0] n750;
  wire [34-1:0] n751;
  wire [34-1:0] n752;
  wire [34-1:0] n753;
  wire [34-1:0] n754;
  wire [34-1:0] n755;
  wire [34-1:0] n756;
  wire [34-1:0] n757;
  wire [34-1:0] n758;
  wire [34-1:0] n759;
  wire [34-1:0] n76;
  wire [34-1:0] n760;
  wire [34-1:0] n761;
  wire [34-1:0] n762;
  wire [34-1:0] n763;
  wire [34-1:0] n764;
  wire [34-1:0] n765;
  wire [34-1:0] n766;
  wire [34-1:0] n767;
  wire [34-1:0] n768;
  wire [34-1:0] n769;
  wire [34-1:0] n77;
  wire [34-1:0] n770;
  wire [34-1:0] n771;
  wire [34-1:0] n772;
  wire [34-1:0] n773;
  wire [34-1:0] n774;
  wire [34-1:0] n775;
  wire [34-1:0] n776;
  wire [34-1:0] n777;
  wire [34-1:0] n778;
  wire [34-1:0] n779;
  wire [34-1:0] n78;
  wire [34-1:0] n780;
  wire [34-1:0] n781;
  wire [34-1:0] n782;
  wire [34-1:0] n783;
  wire [34-1:0] n784;
  wire [34-1:0] n785;
  wire [34-1:0] n786;
  wire [34-1:0] n787;
  wire [34-1:0] n788;
  wire [34-1:0] n789;
  wire [34-1:0] n79;
  wire [34-1:0] n790;
  wire [34-1:0] n791;
  wire [34-1:0] n792;
  wire [34-1:0] n793;
  wire [34-1:0] n794;
  wire [34-1:0] n795;
  wire [34-1:0] n796;
  wire [34-1:0] n797;
  wire [34-1:0] n798;
  wire [34-1:0] n799;
  wire [34-1:0] n8;
  wire [34-1:0] n80;
  wire [34-1:0] n800;
  wire [34-1:0] n801;
  wire [34-1:0] n802;
  wire [34-1:0] n803;
  wire [34-1:0] n804;
  wire [34-1:0] n805;
  wire [34-1:0] n806;
  wire [34-1:0] n807;
  wire [34-1:0] n808;
  wire [34-1:0] n809;
  wire [34-1:0] n81;
  wire [34-1:0] n810;
  wire [34-1:0] n811;
  wire [34-1:0] n812;
  wire [34-1:0] n813;
  wire [34-1:0] n814;
  wire [34-1:0] n815;
  wire [34-1:0] n816;
  wire [34-1:0] n817;
  wire [34-1:0] n818;
  wire [34-1:0] n819;
  wire [34-1:0] n82;
  wire [34-1:0] n820;
  wire [34-1:0] n821;
  wire [34-1:0] n822;
  wire [34-1:0] n823;
  wire [34-1:0] n824;
  wire [34-1:0] n825;
  wire [34-1:0] n826;
  wire [34-1:0] n827;
  wire [34-1:0] n828;
  wire [34-1:0] n829;
  wire [34-1:0] n83;
  wire [34-1:0] n830;
  wire [34-1:0] n831;
  wire [34-1:0] n832;
  wire [34-1:0] n833;
  wire [34-1:0] n834;
  wire [34-1:0] n835;
  wire [34-1:0] n836;
  wire [34-1:0] n837;
  wire [34-1:0] n838;
  wire [34-1:0] n839;
  wire [34-1:0] n84;
  wire [34-1:0] n840;
  wire [34-1:0] n841;
  wire [34-1:0] n842;
  wire [34-1:0] n843;
  wire [34-1:0] n844;
  wire [34-1:0] n845;
  wire [34-1:0] n846;
  wire [34-1:0] n847;
  wire [34-1:0] n848;
  wire [34-1:0] n849;
  wire [34-1:0] n85;
  wire [34-1:0] n850;
  wire [34-1:0] n851;
  wire [34-1:0] n852;
  wire [34-1:0] n853;
  wire [34-1:0] n854;
  wire [34-1:0] n855;
  wire [34-1:0] n856;
  wire [34-1:0] n857;
  wire [34-1:0] n858;
  wire [34-1:0] n859;
  wire [34-1:0] n86;
  wire [34-1:0] n860;
  wire [34-1:0] n861;
  wire [34-1:0] n862;
  wire [34-1:0] n863;
  wire [34-1:0] n864;
  wire [34-1:0] n865;
  wire [34-1:0] n866;
  wire [34-1:0] n867;
  wire [34-1:0] n868;
  wire [34-1:0] n869;
  wire [34-1:0] n87;
  wire [34-1:0] n870;
  wire [34-1:0] n871;
  wire [34-1:0] n872;
  wire [34-1:0] n873;
  wire [34-1:0] n874;
  wire [34-1:0] n875;
  wire [34-1:0] n876;
  wire [34-1:0] n877;
  wire [34-1:0] n878;
  wire [34-1:0] n879;
  wire [34-1:0] n88;
  wire [34-1:0] n880;
  wire [34-1:0] n881;
  wire [34-1:0] n882;
  wire [34-1:0] n883;
  wire [34-1:0] n884;
  wire [34-1:0] n885;
  wire [34-1:0] n886;
  wire [34-1:0] n887;
  wire [34-1:0] n888;
  wire [34-1:0] n889;
  wire [34-1:0] n89;
  wire [34-1:0] n890;
  wire [34-1:0] n891;
  wire [34-1:0] n892;
  wire [34-1:0] n893;
  wire [34-1:0] n894;
  wire [34-1:0] n895;
  wire [34-1:0] n896;
  wire [34-1:0] n897;
  wire [34-1:0] n898;
  wire [34-1:0] n899;
  wire [34-1:0] n9;
  wire [34-1:0] n90;
  wire [34-1:0] n900;
  wire [34-1:0] n901;
  wire [34-1:0] n902;
  wire [34-1:0] n903;
  wire [34-1:0] n904;
  wire [34-1:0] n905;
  wire [34-1:0] n906;
  wire [34-1:0] n907;
  wire [34-1:0] n908;
  wire [34-1:0] n909;
  wire [34-1:0] n91;
  wire [34-1:0] n910;
  wire [34-1:0] n911;
  wire [34-1:0] n912;
  wire [34-1:0] n913;
  wire [34-1:0] n914;
  wire [34-1:0] n915;
  wire [34-1:0] n916;
  wire [34-1:0] n917;
  wire [34-1:0] n918;
  wire [34-1:0] n919;
  wire [34-1:0] n92;
  wire [34-1:0] n920;
  wire [34-1:0] n921;
  wire [34-1:0] n922;
  wire [34-1:0] n923;
  wire [34-1:0] n924;
  wire [34-1:0] n925;
  wire [34-1:0] n926;
  wire [34-1:0] n927;
  wire [34-1:0] n928;
  wire [34-1:0] n929;
  wire [34-1:0] n93;
  wire [34-1:0] n930;
  wire [34-1:0] n931;
  wire [34-1:0] n932;
  wire [34-1:0] n933;
  wire [34-1:0] n934;
  wire [34-1:0] n935;
  wire [34-1:0] n936;
  wire [34-1:0] n937;
  wire [34-1:0] n938;
  wire [34-1:0] n939;
  wire [34-1:0] n94;
  wire [34-1:0] n940;
  wire [34-1:0] n941;
  wire [34-1:0] n942;
  wire [34-1:0] n943;
  wire [34-1:0] n944;
  wire [34-1:0] n945;
  wire [34-1:0] n946;
  wire [34-1:0] n947;
  wire [34-1:0] n948;
  wire [34-1:0] n949;
  wire [34-1:0] n95;
  wire [34-1:0] n950;
  wire [34-1:0] n951;
  wire [34-1:0] n952;
  wire [34-1:0] n953;
  wire [34-1:0] n954;
  wire [34-1:0] n955;
  wire [34-1:0] n956;
  wire [34-1:0] n957;
  wire [34-1:0] n958;
  wire [34-1:0] n959;
  wire [34-1:0] n96;
  wire [34-1:0] n960;
  wire [34-1:0] n961;
  wire [34-1:0] n962;
  wire [34-1:0] n963;
  wire [34-1:0] n964;
  wire [34-1:0] n965;
  wire [34-1:0] n966;
  wire [34-1:0] n967;
  wire [34-1:0] n968;
  wire [34-1:0] n969;
  wire [34-1:0] n97;
  wire [34-1:0] n970;
  wire [34-1:0] n971;
  wire [34-1:0] n972;
  wire [34-1:0] n973;
  wire [34-1:0] n974;
  wire [34-1:0] n975;
  wire [34-1:0] n976;
  wire [34-1:0] n977;
  wire [34-1:0] n978;
  wire [34-1:0] n979;
  wire [34-1:0] n98;
  wire [34-1:0] n980;
  wire [34-1:0] n981;
  wire [34-1:0] n982;
  wire [34-1:0] n983;
  wire [34-1:0] n984;
  wire [34-1:0] n985;
  wire [34-1:0] n986;
  wire [34-1:0] n987;
  wire [34-1:0] n988;
  wire [34-1:0] n989;
  wire [34-1:0] n99;
  wire [34-1:0] n990;
  wire [34-1:0] n991;
  wire [34-1:0] n992;
  wire [34-1:0] n993;
  wire [34-1:0] n994;
  wire [34-1:0] n995;
  wire [34-1:0] n996;
  wire [34-1:0] n997;
  wire [34-1:0] n998;
  wire [34-1:0] n999;
  wire [4-1:0] streams_ready;
  wire en;
  assign en = &streams_ready;
  wire [2-1:0] done_wire;

  always @(posedge clk) begin
    acc_user_done <= &done_wire;
  end


  SyncAdd
  add_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1242),
    .din1(n1265),
    .dout0(n1302)
  );


  SyncAdd
  add_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1241),
    .din1(n1251),
    .dout0(n1252)
  );


  SyncAdd
  add_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1430),
    .din1(n1453),
    .dout0(n1492)
  );


  SyncAdd
  add_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1429),
    .din1(n1439),
    .dout0(n1440)
  );


  SyncAdd
  add_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1468),
    .din1(n1491),
    .dout0(n1530)
  );


  SyncAdd
  add_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1467),
    .din1(n1477),
    .dout0(n1478)
  );


  SyncAdd
  add_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1506),
    .din1(n1529),
    .dout0(n1568)
  );


  SyncAdd
  add_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1505),
    .din1(n1515),
    .dout0(n1516)
  );


  SyncAdd
  add_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1544),
    .din1(n1567),
    .dout0(n1606)
  );


  SyncAdd
  add_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1543),
    .din1(n1553),
    .dout0(n1554)
  );


  SyncAdd
  add_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1582),
    .din1(n1605),
    .dout0(n1644)
  );


  SyncAdd
  add_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1581),
    .din1(n1591),
    .dout0(n1592)
  );


  SyncAdd
  add_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1278),
    .din1(n1301),
    .dout0(n1340)
  );


  SyncAdd
  add_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1620),
    .din1(n1643),
    .dout0(n1682)
  );


  SyncAdd
  add_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1619),
    .din1(n1629),
    .dout0(n1630)
  );


  SyncAdd
  add_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1658),
    .din1(n1681),
    .dout0(n1720)
  );


  SyncAdd
  add_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1657),
    .din1(n1667),
    .dout0(n1668)
  );


  SyncAdd
  add_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1696),
    .din1(n1719),
    .dout0(n1758)
  );


  SyncAdd
  add_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1695),
    .din1(n1705),
    .dout0(n1706)
  );


  SyncAdd
  add_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1734),
    .din1(n1757),
    .dout0(n1796)
  );


  SyncAdd
  add_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1733),
    .din1(n1743),
    .dout0(n1744)
  );


  SyncAdd
  add_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1772),
    .din1(n1795),
    .dout0(n1834)
  );


  SyncAdd
  add_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1771),
    .din1(n1781),
    .dout0(n1782)
  );


  SyncAdd
  add_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1277),
    .din1(n1287),
    .dout0(n1288)
  );


  SyncAdd
  add_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1810),
    .din1(n1833),
    .dout0(n1872)
  );


  SyncAdd
  add_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1809),
    .din1(n1819),
    .dout0(n1820)
  );


  SyncAdd
  add_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1848),
    .din1(n1871),
    .dout0(n1910)
  );


  SyncAdd
  add_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1847),
    .din1(n1857),
    .dout0(n1858)
  );


  SyncAdd
  add_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1886),
    .din1(n1909),
    .dout0(n1948)
  );


  SyncAdd
  add_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1885),
    .din1(n1895),
    .dout0(n1896)
  );


  SyncAdd
  add_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1924),
    .din1(n1947),
    .dout0(n1986)
  );


  SyncAdd
  add_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1923),
    .din1(n1933),
    .dout0(n1934)
  );


  SyncAdd
  add_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1962),
    .din1(n1985),
    .dout0(n2024)
  );


  SyncAdd
  add_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1961),
    .din1(n1971),
    .dout0(n1972)
  );


  SyncAdd
  add_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1316),
    .din1(n1339),
    .dout0(n1378)
  );


  SyncAdd
  add_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2000),
    .din1(n2023),
    .dout0(n2062)
  );


  SyncAdd
  add_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1999),
    .din1(n2009),
    .dout0(n2010)
  );


  SyncAdd
  add_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2038),
    .din1(n2061),
    .dout0(n2100)
  );


  SyncAdd
  add_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2037),
    .din1(n2047),
    .dout0(n2048)
  );


  SyncAdd
  add_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2076),
    .din1(n2099),
    .dout0(n2138)
  );


  SyncAdd
  add_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2075),
    .din1(n2085),
    .dout0(n2086)
  );


  SyncAdd
  add_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2114),
    .din1(n2137),
    .dout0(n2176)
  );


  SyncAdd
  add_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2113),
    .din1(n2123),
    .dout0(n2124)
  );


  SyncAdd
  add_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2152),
    .din1(n2175),
    .dout0(n2214)
  );


  SyncAdd
  add_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2151),
    .din1(n2161),
    .dout0(n2162)
  );


  SyncAdd
  add_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1315),
    .din1(n1325),
    .dout0(n1326)
  );


  SyncAdd
  add_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2190),
    .din1(n2213),
    .dout0(n2252)
  );


  SyncAdd
  add_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2189),
    .din1(n2199),
    .dout0(n2200)
  );


  SyncAdd
  add_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2228),
    .din1(n2251),
    .dout0(n2290)
  );


  SyncAdd
  add_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2227),
    .din1(n2237),
    .dout0(n2238)
  );


  SyncAdd
  add_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2266),
    .din1(n2289),
    .dout0(n2328)
  );


  SyncAdd
  add_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2265),
    .din1(n2275),
    .dout0(n2276)
  );


  SyncAdd
  add_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2304),
    .din1(n2327),
    .dout0(n2366)
  );


  SyncAdd
  add_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2303),
    .din1(n2313),
    .dout0(n2314)
  );


  SyncAdd
  add_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2342),
    .din1(n2365),
    .dout0(n2404)
  );


  SyncAdd
  add_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2341),
    .din1(n2351),
    .dout0(n2352)
  );


  SyncAdd
  add_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1354),
    .din1(n1377),
    .dout0(n1416)
  );


  SyncAdd
  add_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2380),
    .din1(n2403),
    .dout0(n2442)
  );


  SyncAdd
  add_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2379),
    .din1(n2389),
    .dout0(n2390)
  );


  SyncAdd
  add_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2418),
    .din1(n2441),
    .dout0(n2448)
  );


  SyncAdd
  add_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2417),
    .din1(n2427),
    .dout0(n2428)
  );


  SyncAdd
  add_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1353),
    .din1(n1363),
    .dout0(n1364)
  );


  SyncAdd
  add_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1392),
    .din1(n1415),
    .dout0(n1454)
  );


  SyncAdd
  add_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1391),
    .din1(n1401),
    .dout0(n1402)
  );


  SyncAdd
  add_fir0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1218),
    .dout0(n1220),
    .din1(n1224)
  );


  SyncAdd
  add_fir1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1220),
    .dout0(n1221),
    .din1(n1225)
  );


  SyncAdd
  add_fir2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1221),
    .din1(n1226),
    .dout0(n2447)
  );


  SyncAdd
  add_fir3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1219),
    .dout0(n1222),
    .din1(n1227)
  );


  SyncAdd
  add_fir4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1222),
    .dout0(n1223),
    .din1(n1228)
  );


  SyncAdd
  add_fir5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1223),
    .din1(n1229),
    .dout0(n2446)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1243),
    .dout0(n1248)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2654435769)
  )
  addi_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1244),
    .dout0(n1247)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1013904242)
  )
  addi_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1295),
    .dout0(n1298)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2175735113)
  )
  addi_C100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1865),
    .dout0(n1868)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1864),
    .dout0(n1866)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1887),
    .dout0(n1892)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(535203586)
  )
  addi_C103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1888),
    .dout0(n1891)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1889),
    .dout0(n1890)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1901),
    .dout0(n1905)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(535203586)
  )
  addi_C106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1903),
    .dout0(n1906)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1902),
    .dout0(n1904)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1925),
    .dout0(n1930)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3189639355)
  )
  addi_C109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1926),
    .dout0(n1929)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1294),
    .dout0(n1296)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1927),
    .dout0(n1928)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1939),
    .dout0(n1943)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3189639355)
  )
  addi_C112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1941),
    .dout0(n1944)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1940),
    .dout0(n1942)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1963),
    .dout0(n1968)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1549107828)
  )
  addi_C115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1964),
    .dout0(n1967)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1965),
    .dout0(n1966)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1977),
    .dout0(n1981)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1549107828)
  )
  addi_C118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1979),
    .dout0(n1982)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1978),
    .dout0(n1980)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1317),
    .dout0(n1322)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2001),
    .dout0(n2006)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4203543597)
  )
  addi_C121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2002),
    .dout0(n2005)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2003),
    .dout0(n2004)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2015),
    .dout0(n2019)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4203543597)
  )
  addi_C124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2017),
    .dout0(n2020)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2016),
    .dout0(n2018)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2039),
    .dout0(n2044)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2563012070)
  )
  addi_C127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2040),
    .dout0(n2043)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C128
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2041),
    .dout0(n2042)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C129
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2053),
    .dout0(n2057)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3668340011)
  )
  addi_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1318),
    .dout0(n1321)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2563012070)
  )
  addi_C130
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2055),
    .dout0(n2058)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C131
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2054),
    .dout0(n2056)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C132
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2077),
    .dout0(n2082)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(922480543)
  )
  addi_C133
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2078),
    .dout0(n2081)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C134
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2079),
    .dout0(n2080)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C135
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2091),
    .dout0(n2095)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(922480543)
  )
  addi_C136
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2093),
    .dout0(n2096)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C137
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2092),
    .dout0(n2094)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C138
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2115),
    .dout0(n2120)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3576916312)
  )
  addi_C139
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2116),
    .dout0(n2119)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1319),
    .dout0(n1320)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C140
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2117),
    .dout0(n2118)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C141
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2129),
    .dout0(n2133)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3576916312)
  )
  addi_C142
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2131),
    .dout0(n2134)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C143
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2130),
    .dout0(n2132)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C144
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2153),
    .dout0(n2158)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1936384785)
  )
  addi_C145
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2154),
    .dout0(n2157)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C146
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2155),
    .dout0(n2156)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C147
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2167),
    .dout0(n2171)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1936384785)
  )
  addi_C148
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2169),
    .dout0(n2172)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C149
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2168),
    .dout0(n2170)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1331),
    .dout0(n1335)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C150
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2191),
    .dout0(n2196)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(295853258)
  )
  addi_C151
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2192),
    .dout0(n2195)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C152
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2193),
    .dout0(n2194)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C153
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2205),
    .dout0(n2209)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(295853258)
  )
  addi_C154
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2207),
    .dout0(n2210)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C155
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2206),
    .dout0(n2208)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C156
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2229),
    .dout0(n2234)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2950289027)
  )
  addi_C157
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2230),
    .dout0(n2233)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C158
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2231),
    .dout0(n2232)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C159
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2243),
    .dout0(n2247)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3668340011)
  )
  addi_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1333),
    .dout0(n1336)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2950289027)
  )
  addi_C160
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2245),
    .dout0(n2248)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C161
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2244),
    .dout0(n2246)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C162
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2267),
    .dout0(n2272)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1309757500)
  )
  addi_C163
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2268),
    .dout0(n2271)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C164
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2269),
    .dout0(n2270)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C165
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2281),
    .dout0(n2285)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1309757500)
  )
  addi_C166
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2283),
    .dout0(n2286)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C167
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2282),
    .dout0(n2284)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C168
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2305),
    .dout0(n2310)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3964193269)
  )
  addi_C169
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2306),
    .dout0(n2309)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1332),
    .dout0(n1334)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C170
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2307),
    .dout0(n2308)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C171
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2319),
    .dout0(n2323)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3964193269)
  )
  addi_C172
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2321),
    .dout0(n2324)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C173
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2320),
    .dout0(n2322)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C174
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2343),
    .dout0(n2348)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2323661742)
  )
  addi_C175
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2344),
    .dout0(n2347)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C176
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2345),
    .dout0(n2346)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C177
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2357),
    .dout0(n2361)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2323661742)
  )
  addi_C178
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2359),
    .dout0(n2362)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C179
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2358),
    .dout0(n2360)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1355),
    .dout0(n1360)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C180
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2381),
    .dout0(n2386)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(683130215)
  )
  addi_C181
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2382),
    .dout0(n2385)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C182
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2383),
    .dout0(n2384)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C183
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2395),
    .dout0(n2399)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(683130215)
  )
  addi_C184
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2397),
    .dout0(n2400)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C185
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2396),
    .dout0(n2398)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C186
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2419),
    .dout0(n2424)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3337565984)
  )
  addi_C187
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2420),
    .dout0(n2423)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C188
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2421),
    .dout0(n2422)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C189
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2433),
    .dout0(n2437)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2027808484)
  )
  addi_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1356),
    .dout0(n1359)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3337565984)
  )
  addi_C190
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2435),
    .dout0(n2438)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C191
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2434),
    .dout0(n2436)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1245),
    .dout0(n1246)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1357),
    .dout0(n1358)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1369),
    .dout0(n1373)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2027808484)
  )
  addi_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1371),
    .dout0(n1374)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1370),
    .dout0(n1372)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1393),
    .dout0(n1398)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(387276957)
  )
  addi_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1394),
    .dout0(n1397)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1395),
    .dout0(n1396)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1407),
    .dout0(n1411)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(387276957)
  )
  addi_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1409),
    .dout0(n1412)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1408),
    .dout0(n1410)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1257),
    .dout0(n1261)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1431),
    .dout0(n1436)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3041712726)
  )
  addi_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1432),
    .dout0(n1435)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1433),
    .dout0(n1434)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1445),
    .dout0(n1449)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3041712726)
  )
  addi_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1447),
    .dout0(n1450)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1446),
    .dout0(n1448)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1469),
    .dout0(n1474)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1401181199)
  )
  addi_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1470),
    .dout0(n1473)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1471),
    .dout0(n1472)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1483),
    .dout0(n1487)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2654435769)
  )
  addi_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1259),
    .dout0(n1262)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1401181199)
  )
  addi_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1485),
    .dout0(n1488)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1484),
    .dout0(n1486)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1507),
    .dout0(n1512)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4055616968)
  )
  addi_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1508),
    .dout0(n1511)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1509),
    .dout0(n1510)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1521),
    .dout0(n1525)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4055616968)
  )
  addi_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1523),
    .dout0(n1526)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1522),
    .dout0(n1524)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1545),
    .dout0(n1550)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2415085441)
  )
  addi_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1546),
    .dout0(n1549)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1258),
    .dout0(n1260)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1547),
    .dout0(n1548)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1559),
    .dout0(n1563)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2415085441)
  )
  addi_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1561),
    .dout0(n1564)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1560),
    .dout0(n1562)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1583),
    .dout0(n1588)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(774553914)
  )
  addi_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1584),
    .dout0(n1587)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1585),
    .dout0(n1586)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1597),
    .dout0(n1601)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(774553914)
  )
  addi_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1599),
    .dout0(n1602)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1598),
    .dout0(n1600)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1279),
    .dout0(n1284)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1621),
    .dout0(n1626)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3428989683)
  )
  addi_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1622),
    .dout0(n1625)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1623),
    .dout0(n1624)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1635),
    .dout0(n1639)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3428989683)
  )
  addi_C64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1637),
    .dout0(n1640)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1636),
    .dout0(n1638)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1659),
    .dout0(n1664)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1788458156)
  )
  addi_C67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1660),
    .dout0(n1663)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1661),
    .dout0(n1662)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1673),
    .dout0(n1677)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1013904242)
  )
  addi_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1280),
    .dout0(n1283)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1788458156)
  )
  addi_C70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1675),
    .dout0(n1678)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1674),
    .dout0(n1676)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1697),
    .dout0(n1702)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(147926629)
  )
  addi_C73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1698),
    .dout0(n1701)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1699),
    .dout0(n1700)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1711),
    .dout0(n1715)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(147926629)
  )
  addi_C76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1713),
    .dout0(n1716)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1712),
    .dout0(n1714)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1735),
    .dout0(n1740)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2802362398)
  )
  addi_C79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1736),
    .dout0(n1739)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1281),
    .dout0(n1282)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1737),
    .dout0(n1738)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1749),
    .dout0(n1753)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2802362398)
  )
  addi_C82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1751),
    .dout0(n1754)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1750),
    .dout0(n1752)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1773),
    .dout0(n1778)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1161830871)
  )
  addi_C85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1774),
    .dout0(n1777)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1775),
    .dout0(n1776)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1787),
    .dout0(n1791)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1161830871)
  )
  addi_C88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1789),
    .dout0(n1792)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1788),
    .dout0(n1790)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1293),
    .dout0(n1297)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1811),
    .dout0(n1816)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3816266640)
  )
  addi_C91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1812),
    .dout0(n1815)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1813),
    .dout0(n1814)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1825),
    .dout0(n1829)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3816266640)
  )
  addi_C94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1827),
    .dout0(n1830)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_C95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1826),
    .dout0(n1828)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_C96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1849),
    .dout0(n1854)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2175735113)
  )
  addi_C97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1850),
    .dout0(n1853)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_C98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1851),
    .dout0(n1852)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_C99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1863),
    .dout0(n1867)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n13),
    .dout0(n18)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3337565984)
  )
  addi_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n14),
    .dout0(n17)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(683130215)
  )
  addi_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n65),
    .dout0(n68)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3816266640)
  )
  addi_D100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n635),
    .dout0(n638)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n634),
    .dout0(n636)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n657),
    .dout0(n662)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1161830871)
  )
  addi_D103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n658),
    .dout0(n661)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n659),
    .dout0(n660)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n671),
    .dout0(n675)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1161830871)
  )
  addi_D106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n673),
    .dout0(n676)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n672),
    .dout0(n674)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n695),
    .dout0(n700)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2802362398)
  )
  addi_D109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n696),
    .dout0(n699)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n64),
    .dout0(n66)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n697),
    .dout0(n698)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n709),
    .dout0(n713)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2802362398)
  )
  addi_D112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n711),
    .dout0(n714)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n710),
    .dout0(n712)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n733),
    .dout0(n738)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(147926629)
  )
  addi_D115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n734),
    .dout0(n737)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n735),
    .dout0(n736)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n747),
    .dout0(n751)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(147926629)
  )
  addi_D118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n749),
    .dout0(n752)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n748),
    .dout0(n750)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n87),
    .dout0(n92)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n771),
    .dout0(n776)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1788458156)
  )
  addi_D121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n772),
    .dout0(n775)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n773),
    .dout0(n774)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n785),
    .dout0(n789)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1788458156)
  )
  addi_D124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n787),
    .dout0(n790)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n786),
    .dout0(n788)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n809),
    .dout0(n814)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3428989683)
  )
  addi_D127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n810),
    .dout0(n813)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D128
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n811),
    .dout0(n812)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D129
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n823),
    .dout0(n827)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2323661742)
  )
  addi_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n88),
    .dout0(n91)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3428989683)
  )
  addi_D130
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n825),
    .dout0(n828)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D131
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n824),
    .dout0(n826)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D132
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n847),
    .dout0(n852)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(774553914)
  )
  addi_D133
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n848),
    .dout0(n851)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D134
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n849),
    .dout0(n850)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D135
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n861),
    .dout0(n865)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(774553914)
  )
  addi_D136
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n863),
    .dout0(n866)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D137
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n862),
    .dout0(n864)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D138
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n885),
    .dout0(n890)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2415085441)
  )
  addi_D139
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n886),
    .dout0(n889)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n89),
    .dout0(n90)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D140
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n887),
    .dout0(n888)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D141
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n899),
    .dout0(n903)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2415085441)
  )
  addi_D142
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n901),
    .dout0(n904)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D143
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n900),
    .dout0(n902)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D144
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n923),
    .dout0(n928)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4055616968)
  )
  addi_D145
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n924),
    .dout0(n927)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D146
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n925),
    .dout0(n926)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D147
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n937),
    .dout0(n941)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4055616968)
  )
  addi_D148
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n939),
    .dout0(n942)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D149
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n938),
    .dout0(n940)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n101),
    .dout0(n105)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D150
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n961),
    .dout0(n966)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1401181199)
  )
  addi_D151
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n962),
    .dout0(n965)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D152
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n963),
    .dout0(n964)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D153
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n975),
    .dout0(n979)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1401181199)
  )
  addi_D154
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n977),
    .dout0(n980)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D155
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n976),
    .dout0(n978)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D156
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1004),
    .din0(n999)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3041712726)
  )
  addi_D157
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1000),
    .dout0(n1003)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D158
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1001),
    .dout0(n1002)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D159
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1013),
    .dout0(n1017)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2323661742)
  )
  addi_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n103),
    .dout0(n106)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3041712726)
  )
  addi_D160
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1015),
    .dout0(n1018)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D161
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1014),
    .dout0(n1016)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D162
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1037),
    .dout0(n1042)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(387276957)
  )
  addi_D163
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1038),
    .dout0(n1041)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D164
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1039),
    .dout0(n1040)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D165
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1051),
    .dout0(n1055)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(387276957)
  )
  addi_D166
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1053),
    .dout0(n1056)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D167
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1052),
    .dout0(n1054)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D168
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1075),
    .dout0(n1080)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2027808484)
  )
  addi_D169
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1076),
    .dout0(n1079)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n102),
    .dout0(n104)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D170
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1077),
    .dout0(n1078)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D171
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1089),
    .dout0(n1093)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2027808484)
  )
  addi_D172
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1091),
    .dout0(n1094)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D173
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1090),
    .dout0(n1092)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D174
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1113),
    .dout0(n1118)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3668340011)
  )
  addi_D175
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1114),
    .dout0(n1117)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D176
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1115),
    .dout0(n1116)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D177
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1127),
    .dout0(n1131)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3668340011)
  )
  addi_D178
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1129),
    .dout0(n1132)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D179
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1128),
    .dout0(n1130)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n125),
    .dout0(n130)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D180
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1151),
    .dout0(n1156)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1013904242)
  )
  addi_D181
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1152),
    .dout0(n1155)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D182
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1153),
    .dout0(n1154)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D183
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1165),
    .dout0(n1169)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1013904242)
  )
  addi_D184
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1167),
    .dout0(n1170)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D185
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1166),
    .dout0(n1168)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D186
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1189),
    .dout0(n1194)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2654435769)
  )
  addi_D187
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1190),
    .dout0(n1193)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D188
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1191),
    .dout0(n1192)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D189
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1203),
    .dout0(n1207)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3964193269)
  )
  addi_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n126),
    .dout0(n129)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2654435769)
  )
  addi_D190
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1205),
    .dout0(n1208)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D191
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1204),
    .dout0(n1206)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n15),
    .dout0(n16)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n127),
    .dout0(n128)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n139),
    .dout0(n143)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3964193269)
  )
  addi_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n141),
    .dout0(n144)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n140),
    .dout0(n142)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n163),
    .dout0(n168)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1309757500)
  )
  addi_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n164),
    .dout0(n167)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n165),
    .dout0(n166)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n177),
    .dout0(n181)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1309757500)
  )
  addi_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n179),
    .dout0(n182)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n178),
    .dout0(n180)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n27),
    .dout0(n31)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n201),
    .dout0(n206)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2950289027)
  )
  addi_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n202),
    .dout0(n205)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n203),
    .dout0(n204)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n215),
    .dout0(n219)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2950289027)
  )
  addi_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n217),
    .dout0(n220)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n216),
    .dout0(n218)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n239),
    .dout0(n244)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(295853258)
  )
  addi_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n240),
    .dout0(n243)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n241),
    .dout0(n242)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n253),
    .dout0(n257)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3337565984)
  )
  addi_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n29),
    .dout0(n32)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(295853258)
  )
  addi_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n255),
    .dout0(n258)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n254),
    .dout0(n256)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n277),
    .dout0(n282)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1936384785)
  )
  addi_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n278),
    .dout0(n281)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n279),
    .dout0(n280)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n291),
    .dout0(n295)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1936384785)
  )
  addi_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n293),
    .dout0(n296)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n292),
    .dout0(n294)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n315),
    .dout0(n320)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3576916312)
  )
  addi_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n316),
    .dout0(n319)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n28),
    .dout0(n30)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n317),
    .dout0(n318)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n329),
    .dout0(n333)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3576916312)
  )
  addi_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n331),
    .dout0(n334)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n330),
    .dout0(n332)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n353),
    .dout0(n358)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(922480543)
  )
  addi_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n354),
    .dout0(n357)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n355),
    .dout0(n356)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n367),
    .dout0(n371)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(922480543)
  )
  addi_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n369),
    .dout0(n372)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n368),
    .dout0(n370)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n49),
    .dout0(n54)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n391),
    .dout0(n396)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2563012070)
  )
  addi_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n392),
    .dout0(n395)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n393),
    .dout0(n394)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n405),
    .dout0(n409)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2563012070)
  )
  addi_D64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n407),
    .dout0(n410)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n406),
    .dout0(n408)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n429),
    .dout0(n434)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4203543597)
  )
  addi_D67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n430),
    .dout0(n433)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n431),
    .dout0(n432)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n443),
    .dout0(n447)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(683130215)
  )
  addi_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n50),
    .dout0(n53)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4203543597)
  )
  addi_D70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n445),
    .dout0(n448)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n444),
    .dout0(n446)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n467),
    .dout0(n472)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1549107828)
  )
  addi_D73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n468),
    .dout0(n471)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n469),
    .dout0(n470)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n481),
    .dout0(n485)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1549107828)
  )
  addi_D76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n483),
    .dout0(n486)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n482),
    .dout0(n484)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n505),
    .dout0(n510)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3189639355)
  )
  addi_D79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n506),
    .dout0(n509)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n51),
    .dout0(n52)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n507),
    .dout0(n508)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n519),
    .dout0(n523)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3189639355)
  )
  addi_D82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n521),
    .dout0(n524)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n520),
    .dout0(n522)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n543),
    .dout0(n548)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(535203586)
  )
  addi_D85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n544),
    .dout0(n547)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n545),
    .dout0(n546)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n557),
    .dout0(n561)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(535203586)
  )
  addi_D88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n559),
    .dout0(n562)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n558),
    .dout0(n560)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n63),
    .dout0(n67)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n581),
    .dout0(n586)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2175735113)
  )
  addi_D91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n582),
    .dout0(n585)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n583),
    .dout0(n584)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n595),
    .dout0(n599)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2175735113)
  )
  addi_D94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n597),
    .dout0(n600)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3342584445)
  )
  addi_D95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n596),
    .dout0(n598)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(1394839874)
  )
  addi_D96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n619),
    .dout0(n624)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(3816266640)
  )
  addi_D97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n620),
    .dout0(n623)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(4089647642)
  )
  addi_D98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n621),
    .dout0(n622)
  );


  SyncAddI
  #(
    .ID(1),
    .IMMEDIATE(2490677480)
  )
  addi_D99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n633),
    .dout0(n637)
  );


  SyncIn
  in0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .start(start),
    .rd_done(acc_user_done_rd_data[0]),
    .rd_available(acc_user_available_read[0]),
    .rd_valid(acc_user_read_data_valid[0]),
    .rd_data(acc_user_read_data[511:0]),
    .rd_en(acc_user_request_read[0]),
    .component_ready(streams_ready[0]),
    .dout0(n2444)
  );


  SyncIn
  in1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .start(start),
    .rd_done(acc_user_done_rd_data[1]),
    .rd_available(acc_user_available_read[1]),
    .rd_valid(acc_user_read_data_valid[1]),
    .rd_data(acc_user_read_data[1023:512]),
    .rd_en(acc_user_request_read[1]),
    .component_ready(streams_ready[1]),
    .dout0(n2445)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(1)
  )
  mult_fir0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1214),
    .dout0(n1216)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  mult_fir1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1214),
    .dout0(n1224)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(3)
  )
  mult_fir2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1214),
    .dout0(n1225)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  mult_fir3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1214),
    .dout0(n1226)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(1)
  )
  mult_fir4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1215),
    .dout0(n1217)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(2)
  )
  mult_fir5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1215),
    .dout0(n1227)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(3)
  )
  mult_fir6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1215),
    .dout0(n1228)
  );


  SyncMulI
  #(
    .ID(1),
    .IMMEDIATE(1)
  )
  mult_fir7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1215),
    .dout0(n1229)
  );


  SyncOut
  out0
  (
    .clk(clk),
    .rst(rst),
    .start(start),
    .en(en),
    .wr_available(acc_user_available_write[0]),
    .wr_data(acc_user_write_data[511:0]),
    .wr_en(acc_user_request_write[0]),
    .component_ready(streams_ready[2]),
    .done(done_wire[0]),
    .din0(n2449)
  );


  SyncOut
  out1
  (
    .clk(clk),
    .rst(rst),
    .start(start),
    .en(en),
    .wr_available(acc_user_available_write[1]),
    .wr_data(acc_user_write_data[1023:512]),
    .wr_en(acc_user_request_write[1]),
    .component_ready(streams_ready[3]),
    .done(done_wire[1]),
    .din0(n2448)
  );


  SyncRegister
  reg_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1230),
    .din0(n2446)
  );


  SyncRegister
  reg_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1238),
    .din0(n2447)
  );


  SyncRegister
  reg_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1234),
    .dout0(n1235)
  );


  SyncRegister
  reg_C100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1402),
    .dout0(n1409)
  );


  SyncRegister
  reg_C101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1385),
    .dout0(n1386)
  );


  SyncRegister
  reg_C102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1403),
    .dout0(n1404)
  );


  SyncRegister
  reg_C103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1386),
    .dout0(n1387)
  );


  SyncRegister
  reg_C104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1404),
    .dout0(n1405)
  );


  SyncRegister
  reg_C105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1387),
    .dout0(n1392)
  );


  SyncRegister
  reg_C106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1405),
    .dout0(n1406)
  );


  SyncRegister
  reg_C107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1406),
    .dout0(n1455)
  );


  SyncRegister
  reg_C108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1396),
    .dout0(n1399)
  );


  SyncRegister
  reg_C109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1410),
    .dout0(n1414)
  );


  SyncRegister
  reg_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1252),
    .dout0(n1253)
  );


  SyncRegister
  reg_C110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1418),
    .din0(n1454)
  );


  SyncRegister
  reg_C111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1426),
    .din0(n1455)
  );


  SyncRegister
  reg_C112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1432),
    .din0(n1454)
  );


  SyncRegister
  reg_C113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1426),
    .dout0(n1427)
  );


  SyncRegister
  reg_C114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1418),
    .dout0(n1419)
  );


  SyncRegister
  reg_C115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1419),
    .dout0(n1420)
  );


  SyncRegister
  reg_C116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1427),
    .dout0(n1428)
  );


  SyncRegister
  reg_C117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1420),
    .dout0(n1421)
  );


  SyncRegister
  reg_C118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1428),
    .dout0(n1429)
  );


  SyncRegister
  reg_C119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1421),
    .dout0(n1422)
  );


  SyncRegister
  reg_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1252),
    .dout0(n1259)
  );


  SyncRegister
  reg_C120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1422),
    .dout0(n1423)
  );


  SyncRegister
  reg_C121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1440),
    .dout0(n1441)
  );


  SyncRegister
  reg_C122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1440),
    .dout0(n1447)
  );


  SyncRegister
  reg_C123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1423),
    .dout0(n1424)
  );


  SyncRegister
  reg_C124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1441),
    .dout0(n1442)
  );


  SyncRegister
  reg_C125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1424),
    .dout0(n1425)
  );


  SyncRegister
  reg_C126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1442),
    .dout0(n1443)
  );


  SyncRegister
  reg_C127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1425),
    .dout0(n1430)
  );


  SyncRegister
  reg_C128
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1443),
    .dout0(n1444)
  );


  SyncRegister
  reg_C129
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1444),
    .dout0(n1493)
  );


  SyncRegister
  reg_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1235),
    .dout0(n1236)
  );


  SyncRegister
  reg_C130
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1434),
    .dout0(n1437)
  );


  SyncRegister
  reg_C131
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1448),
    .dout0(n1452)
  );


  SyncRegister
  reg_C132
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1456),
    .din0(n1492)
  );


  SyncRegister
  reg_C133
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1464),
    .din0(n1493)
  );


  SyncRegister
  reg_C134
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1470),
    .din0(n1492)
  );


  SyncRegister
  reg_C135
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1464),
    .dout0(n1465)
  );


  SyncRegister
  reg_C136
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1456),
    .dout0(n1457)
  );


  SyncRegister
  reg_C137
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1457),
    .dout0(n1458)
  );


  SyncRegister
  reg_C138
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1465),
    .dout0(n1466)
  );


  SyncRegister
  reg_C139
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1458),
    .dout0(n1459)
  );


  SyncRegister
  reg_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1253),
    .dout0(n1254)
  );


  SyncRegister
  reg_C140
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1466),
    .dout0(n1467)
  );


  SyncRegister
  reg_C141
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1459),
    .dout0(n1460)
  );


  SyncRegister
  reg_C142
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1460),
    .dout0(n1461)
  );


  SyncRegister
  reg_C143
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1478),
    .dout0(n1479)
  );


  SyncRegister
  reg_C144
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1478),
    .dout0(n1485)
  );


  SyncRegister
  reg_C145
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1461),
    .dout0(n1462)
  );


  SyncRegister
  reg_C146
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1479),
    .dout0(n1480)
  );


  SyncRegister
  reg_C147
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1462),
    .dout0(n1463)
  );


  SyncRegister
  reg_C148
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1480),
    .dout0(n1481)
  );


  SyncRegister
  reg_C149
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1463),
    .dout0(n1468)
  );


  SyncRegister
  reg_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1236),
    .dout0(n1237)
  );


  SyncRegister
  reg_C150
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1481),
    .dout0(n1482)
  );


  SyncRegister
  reg_C151
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1482),
    .dout0(n1531)
  );


  SyncRegister
  reg_C152
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1472),
    .dout0(n1475)
  );


  SyncRegister
  reg_C153
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1486),
    .dout0(n1490)
  );


  SyncRegister
  reg_C154
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1494),
    .din0(n1530)
  );


  SyncRegister
  reg_C155
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1502),
    .din0(n1531)
  );


  SyncRegister
  reg_C156
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1508),
    .din0(n1530)
  );


  SyncRegister
  reg_C157
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1502),
    .dout0(n1503)
  );


  SyncRegister
  reg_C158
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1494),
    .dout0(n1495)
  );


  SyncRegister
  reg_C159
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1495),
    .dout0(n1496)
  );


  SyncRegister
  reg_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1254),
    .dout0(n1255)
  );


  SyncRegister
  reg_C160
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1503),
    .dout0(n1504)
  );


  SyncRegister
  reg_C161
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1496),
    .dout0(n1497)
  );


  SyncRegister
  reg_C162
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1504),
    .dout0(n1505)
  );


  SyncRegister
  reg_C163
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1497),
    .dout0(n1498)
  );


  SyncRegister
  reg_C164
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1498),
    .dout0(n1499)
  );


  SyncRegister
  reg_C165
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1516),
    .dout0(n1517)
  );


  SyncRegister
  reg_C166
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1516),
    .dout0(n1523)
  );


  SyncRegister
  reg_C167
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1499),
    .dout0(n1500)
  );


  SyncRegister
  reg_C168
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1517),
    .dout0(n1518)
  );


  SyncRegister
  reg_C169
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1500),
    .dout0(n1501)
  );


  SyncRegister
  reg_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1237),
    .dout0(n1242)
  );


  SyncRegister
  reg_C170
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1518),
    .dout0(n1519)
  );


  SyncRegister
  reg_C171
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1501),
    .dout0(n1506)
  );


  SyncRegister
  reg_C172
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1519),
    .dout0(n1520)
  );


  SyncRegister
  reg_C173
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1520),
    .dout0(n1569)
  );


  SyncRegister
  reg_C174
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1510),
    .dout0(n1513)
  );


  SyncRegister
  reg_C175
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1524),
    .dout0(n1528)
  );


  SyncRegister
  reg_C176
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1532),
    .din0(n1568)
  );


  SyncRegister
  reg_C177
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1540),
    .din0(n1569)
  );


  SyncRegister
  reg_C178
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1546),
    .din0(n1568)
  );


  SyncRegister
  reg_C179
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1540),
    .dout0(n1541)
  );


  SyncRegister
  reg_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1255),
    .dout0(n1256)
  );


  SyncRegister
  reg_C180
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1532),
    .dout0(n1533)
  );


  SyncRegister
  reg_C181
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1533),
    .dout0(n1534)
  );


  SyncRegister
  reg_C182
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1541),
    .dout0(n1542)
  );


  SyncRegister
  reg_C183
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1534),
    .dout0(n1535)
  );


  SyncRegister
  reg_C184
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1542),
    .dout0(n1543)
  );


  SyncRegister
  reg_C185
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1535),
    .dout0(n1536)
  );


  SyncRegister
  reg_C186
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1536),
    .dout0(n1537)
  );


  SyncRegister
  reg_C187
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1554),
    .dout0(n1555)
  );


  SyncRegister
  reg_C188
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1554),
    .dout0(n1561)
  );


  SyncRegister
  reg_C189
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1537),
    .dout0(n1538)
  );


  SyncRegister
  reg_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1256),
    .dout0(n1303)
  );


  SyncRegister
  reg_C190
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1555),
    .dout0(n1556)
  );


  SyncRegister
  reg_C191
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1538),
    .dout0(n1539)
  );


  SyncRegister
  reg_C192
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1556),
    .dout0(n1557)
  );


  SyncRegister
  reg_C193
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1539),
    .dout0(n1544)
  );


  SyncRegister
  reg_C194
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1557),
    .dout0(n1558)
  );


  SyncRegister
  reg_C195
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1558),
    .dout0(n1607)
  );


  SyncRegister
  reg_C196
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1548),
    .dout0(n1551)
  );


  SyncRegister
  reg_C197
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1562),
    .dout0(n1566)
  );


  SyncRegister
  reg_C198
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1570),
    .din0(n1606)
  );


  SyncRegister
  reg_C199
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1578),
    .din0(n1607)
  );


  SyncRegister
  reg_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1244),
    .din0(n2446)
  );


  SyncRegister
  reg_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1246),
    .dout0(n1249)
  );


  SyncRegister
  reg_C200
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1584),
    .din0(n1606)
  );


  SyncRegister
  reg_C201
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1578),
    .dout0(n1579)
  );


  SyncRegister
  reg_C202
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1570),
    .dout0(n1571)
  );


  SyncRegister
  reg_C203
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1571),
    .dout0(n1572)
  );


  SyncRegister
  reg_C204
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1579),
    .dout0(n1580)
  );


  SyncRegister
  reg_C205
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1572),
    .dout0(n1573)
  );


  SyncRegister
  reg_C206
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1580),
    .dout0(n1581)
  );


  SyncRegister
  reg_C207
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1573),
    .dout0(n1574)
  );


  SyncRegister
  reg_C208
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1574),
    .dout0(n1575)
  );


  SyncRegister
  reg_C209
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1592),
    .dout0(n1593)
  );


  SyncRegister
  reg_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1260),
    .dout0(n1264)
  );


  SyncRegister
  reg_C210
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1592),
    .dout0(n1599)
  );


  SyncRegister
  reg_C211
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1575),
    .dout0(n1576)
  );


  SyncRegister
  reg_C212
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1593),
    .dout0(n1594)
  );


  SyncRegister
  reg_C213
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1576),
    .dout0(n1577)
  );


  SyncRegister
  reg_C214
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1594),
    .dout0(n1595)
  );


  SyncRegister
  reg_C215
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1577),
    .dout0(n1582)
  );


  SyncRegister
  reg_C216
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1595),
    .dout0(n1596)
  );


  SyncRegister
  reg_C217
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1596),
    .dout0(n1645)
  );


  SyncRegister
  reg_C218
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1586),
    .dout0(n1589)
  );


  SyncRegister
  reg_C219
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1600),
    .dout0(n1604)
  );


  SyncRegister
  reg_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1266),
    .din0(n1302)
  );


  SyncRegister
  reg_C220
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1608),
    .din0(n1644)
  );


  SyncRegister
  reg_C221
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1616),
    .din0(n1645)
  );


  SyncRegister
  reg_C222
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1622),
    .din0(n1644)
  );


  SyncRegister
  reg_C223
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1616),
    .dout0(n1617)
  );


  SyncRegister
  reg_C224
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1608),
    .dout0(n1609)
  );


  SyncRegister
  reg_C225
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1609),
    .dout0(n1610)
  );


  SyncRegister
  reg_C226
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1617),
    .dout0(n1618)
  );


  SyncRegister
  reg_C227
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1610),
    .dout0(n1611)
  );


  SyncRegister
  reg_C228
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1618),
    .dout0(n1619)
  );


  SyncRegister
  reg_C229
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1611),
    .dout0(n1612)
  );


  SyncRegister
  reg_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1274),
    .din0(n1303)
  );


  SyncRegister
  reg_C230
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1612),
    .dout0(n1613)
  );


  SyncRegister
  reg_C231
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1630),
    .dout0(n1631)
  );


  SyncRegister
  reg_C232
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1630),
    .dout0(n1637)
  );


  SyncRegister
  reg_C233
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1613),
    .dout0(n1614)
  );


  SyncRegister
  reg_C234
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1631),
    .dout0(n1632)
  );


  SyncRegister
  reg_C235
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1614),
    .dout0(n1615)
  );


  SyncRegister
  reg_C236
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1632),
    .dout0(n1633)
  );


  SyncRegister
  reg_C237
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1615),
    .dout0(n1620)
  );


  SyncRegister
  reg_C238
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1633),
    .dout0(n1634)
  );


  SyncRegister
  reg_C239
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1634),
    .dout0(n1683)
  );


  SyncRegister
  reg_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1280),
    .din0(n1302)
  );


  SyncRegister
  reg_C240
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1624),
    .dout0(n1627)
  );


  SyncRegister
  reg_C241
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1638),
    .dout0(n1642)
  );


  SyncRegister
  reg_C242
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1646),
    .din0(n1682)
  );


  SyncRegister
  reg_C243
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1654),
    .din0(n1683)
  );


  SyncRegister
  reg_C244
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1660),
    .din0(n1682)
  );


  SyncRegister
  reg_C245
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1654),
    .dout0(n1655)
  );


  SyncRegister
  reg_C246
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1646),
    .dout0(n1647)
  );


  SyncRegister
  reg_C247
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1647),
    .dout0(n1648)
  );


  SyncRegister
  reg_C248
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1655),
    .dout0(n1656)
  );


  SyncRegister
  reg_C249
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1648),
    .dout0(n1649)
  );


  SyncRegister
  reg_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1274),
    .dout0(n1275)
  );


  SyncRegister
  reg_C250
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1656),
    .dout0(n1657)
  );


  SyncRegister
  reg_C251
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1649),
    .dout0(n1650)
  );


  SyncRegister
  reg_C252
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1650),
    .dout0(n1651)
  );


  SyncRegister
  reg_C253
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1668),
    .dout0(n1669)
  );


  SyncRegister
  reg_C254
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1668),
    .dout0(n1675)
  );


  SyncRegister
  reg_C255
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1651),
    .dout0(n1652)
  );


  SyncRegister
  reg_C256
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1669),
    .dout0(n1670)
  );


  SyncRegister
  reg_C257
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1652),
    .dout0(n1653)
  );


  SyncRegister
  reg_C258
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1670),
    .dout0(n1671)
  );


  SyncRegister
  reg_C259
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1653),
    .dout0(n1658)
  );


  SyncRegister
  reg_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1266),
    .dout0(n1267)
  );


  SyncRegister
  reg_C260
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1671),
    .dout0(n1672)
  );


  SyncRegister
  reg_C261
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1672),
    .dout0(n1721)
  );


  SyncRegister
  reg_C262
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1662),
    .dout0(n1665)
  );


  SyncRegister
  reg_C263
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1676),
    .dout0(n1680)
  );


  SyncRegister
  reg_C264
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1684),
    .din0(n1720)
  );


  SyncRegister
  reg_C265
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1692),
    .din0(n1721)
  );


  SyncRegister
  reg_C266
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1698),
    .din0(n1720)
  );


  SyncRegister
  reg_C267
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1692),
    .dout0(n1693)
  );


  SyncRegister
  reg_C268
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1684),
    .dout0(n1685)
  );


  SyncRegister
  reg_C269
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1685),
    .dout0(n1686)
  );


  SyncRegister
  reg_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1267),
    .dout0(n1268)
  );


  SyncRegister
  reg_C270
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1693),
    .dout0(n1694)
  );


  SyncRegister
  reg_C271
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1686),
    .dout0(n1687)
  );


  SyncRegister
  reg_C272
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1694),
    .dout0(n1695)
  );


  SyncRegister
  reg_C273
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1687),
    .dout0(n1688)
  );


  SyncRegister
  reg_C274
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1688),
    .dout0(n1689)
  );


  SyncRegister
  reg_C275
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1706),
    .dout0(n1707)
  );


  SyncRegister
  reg_C276
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1706),
    .dout0(n1713)
  );


  SyncRegister
  reg_C277
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1689),
    .dout0(n1690)
  );


  SyncRegister
  reg_C278
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1707),
    .dout0(n1708)
  );


  SyncRegister
  reg_C279
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1690),
    .dout0(n1691)
  );


  SyncRegister
  reg_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1275),
    .dout0(n1276)
  );


  SyncRegister
  reg_C280
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1708),
    .dout0(n1709)
  );


  SyncRegister
  reg_C281
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1691),
    .dout0(n1696)
  );


  SyncRegister
  reg_C282
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1709),
    .dout0(n1710)
  );


  SyncRegister
  reg_C283
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1710),
    .dout0(n1759)
  );


  SyncRegister
  reg_C284
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1700),
    .dout0(n1703)
  );


  SyncRegister
  reg_C285
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1714),
    .dout0(n1718)
  );


  SyncRegister
  reg_C286
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1722),
    .din0(n1758)
  );


  SyncRegister
  reg_C287
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1730),
    .din0(n1759)
  );


  SyncRegister
  reg_C288
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1736),
    .din0(n1758)
  );


  SyncRegister
  reg_C289
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1730),
    .dout0(n1731)
  );


  SyncRegister
  reg_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1268),
    .dout0(n1269)
  );


  SyncRegister
  reg_C290
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1722),
    .dout0(n1723)
  );


  SyncRegister
  reg_C291
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1723),
    .dout0(n1724)
  );


  SyncRegister
  reg_C292
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1731),
    .dout0(n1732)
  );


  SyncRegister
  reg_C293
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1724),
    .dout0(n1725)
  );


  SyncRegister
  reg_C294
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1732),
    .dout0(n1733)
  );


  SyncRegister
  reg_C295
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1725),
    .dout0(n1726)
  );


  SyncRegister
  reg_C296
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1726),
    .dout0(n1727)
  );


  SyncRegister
  reg_C297
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1744),
    .dout0(n1745)
  );


  SyncRegister
  reg_C298
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1744),
    .dout0(n1751)
  );


  SyncRegister
  reg_C299
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1727),
    .dout0(n1728)
  );


  SyncRegister
  reg_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1238),
    .dout0(n1239)
  );


  SyncRegister
  reg_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1276),
    .dout0(n1277)
  );


  SyncRegister
  reg_C300
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1745),
    .dout0(n1746)
  );


  SyncRegister
  reg_C301
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1728),
    .dout0(n1729)
  );


  SyncRegister
  reg_C302
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1746),
    .dout0(n1747)
  );


  SyncRegister
  reg_C303
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1729),
    .dout0(n1734)
  );


  SyncRegister
  reg_C304
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1747),
    .dout0(n1748)
  );


  SyncRegister
  reg_C305
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1748),
    .dout0(n1797)
  );


  SyncRegister
  reg_C306
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1738),
    .dout0(n1741)
  );


  SyncRegister
  reg_C307
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1752),
    .dout0(n1756)
  );


  SyncRegister
  reg_C308
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1760),
    .din0(n1796)
  );


  SyncRegister
  reg_C309
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1768),
    .din0(n1797)
  );


  SyncRegister
  reg_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1269),
    .dout0(n1270)
  );


  SyncRegister
  reg_C310
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1774),
    .din0(n1796)
  );


  SyncRegister
  reg_C311
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1768),
    .dout0(n1769)
  );


  SyncRegister
  reg_C312
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1760),
    .dout0(n1761)
  );


  SyncRegister
  reg_C313
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1761),
    .dout0(n1762)
  );


  SyncRegister
  reg_C314
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1769),
    .dout0(n1770)
  );


  SyncRegister
  reg_C315
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1762),
    .dout0(n1763)
  );


  SyncRegister
  reg_C316
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1770),
    .dout0(n1771)
  );


  SyncRegister
  reg_C317
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1763),
    .dout0(n1764)
  );


  SyncRegister
  reg_C318
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1764),
    .dout0(n1765)
  );


  SyncRegister
  reg_C319
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1782),
    .dout0(n1783)
  );


  SyncRegister
  reg_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1270),
    .dout0(n1271)
  );


  SyncRegister
  reg_C320
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1782),
    .dout0(n1789)
  );


  SyncRegister
  reg_C321
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1765),
    .dout0(n1766)
  );


  SyncRegister
  reg_C322
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1783),
    .dout0(n1784)
  );


  SyncRegister
  reg_C323
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1766),
    .dout0(n1767)
  );


  SyncRegister
  reg_C324
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1784),
    .dout0(n1785)
  );


  SyncRegister
  reg_C325
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1767),
    .dout0(n1772)
  );


  SyncRegister
  reg_C326
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1785),
    .dout0(n1786)
  );


  SyncRegister
  reg_C327
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1786),
    .dout0(n1835)
  );


  SyncRegister
  reg_C328
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1776),
    .dout0(n1779)
  );


  SyncRegister
  reg_C329
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1790),
    .dout0(n1794)
  );


  SyncRegister
  reg_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1288),
    .dout0(n1289)
  );


  SyncRegister
  reg_C330
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1798),
    .din0(n1834)
  );


  SyncRegister
  reg_C331
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1806),
    .din0(n1835)
  );


  SyncRegister
  reg_C332
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1812),
    .din0(n1834)
  );


  SyncRegister
  reg_C333
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1806),
    .dout0(n1807)
  );


  SyncRegister
  reg_C334
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1798),
    .dout0(n1799)
  );


  SyncRegister
  reg_C335
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1799),
    .dout0(n1800)
  );


  SyncRegister
  reg_C336
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1807),
    .dout0(n1808)
  );


  SyncRegister
  reg_C337
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1800),
    .dout0(n1801)
  );


  SyncRegister
  reg_C338
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1808),
    .dout0(n1809)
  );


  SyncRegister
  reg_C339
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1801),
    .dout0(n1802)
  );


  SyncRegister
  reg_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1288),
    .dout0(n1295)
  );


  SyncRegister
  reg_C340
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1802),
    .dout0(n1803)
  );


  SyncRegister
  reg_C341
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1820),
    .dout0(n1821)
  );


  SyncRegister
  reg_C342
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1820),
    .dout0(n1827)
  );


  SyncRegister
  reg_C343
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1803),
    .dout0(n1804)
  );


  SyncRegister
  reg_C344
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1821),
    .dout0(n1822)
  );


  SyncRegister
  reg_C345
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1804),
    .dout0(n1805)
  );


  SyncRegister
  reg_C346
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1822),
    .dout0(n1823)
  );


  SyncRegister
  reg_C347
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1805),
    .dout0(n1810)
  );


  SyncRegister
  reg_C348
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1823),
    .dout0(n1824)
  );


  SyncRegister
  reg_C349
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1824),
    .dout0(n1873)
  );


  SyncRegister
  reg_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1271),
    .dout0(n1272)
  );


  SyncRegister
  reg_C350
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1814),
    .dout0(n1817)
  );


  SyncRegister
  reg_C351
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1828),
    .dout0(n1832)
  );


  SyncRegister
  reg_C352
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1836),
    .din0(n1872)
  );


  SyncRegister
  reg_C353
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1844),
    .din0(n1873)
  );


  SyncRegister
  reg_C354
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1850),
    .din0(n1872)
  );


  SyncRegister
  reg_C355
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1844),
    .dout0(n1845)
  );


  SyncRegister
  reg_C356
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1836),
    .dout0(n1837)
  );


  SyncRegister
  reg_C357
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1837),
    .dout0(n1838)
  );


  SyncRegister
  reg_C358
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1845),
    .dout0(n1846)
  );


  SyncRegister
  reg_C359
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1838),
    .dout0(n1839)
  );


  SyncRegister
  reg_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1289),
    .dout0(n1290)
  );


  SyncRegister
  reg_C360
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1846),
    .dout0(n1847)
  );


  SyncRegister
  reg_C361
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1839),
    .dout0(n1840)
  );


  SyncRegister
  reg_C362
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1840),
    .dout0(n1841)
  );


  SyncRegister
  reg_C363
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1858),
    .dout0(n1859)
  );


  SyncRegister
  reg_C364
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1858),
    .dout0(n1865)
  );


  SyncRegister
  reg_C365
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1841),
    .dout0(n1842)
  );


  SyncRegister
  reg_C366
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1859),
    .dout0(n1860)
  );


  SyncRegister
  reg_C367
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1842),
    .dout0(n1843)
  );


  SyncRegister
  reg_C368
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1860),
    .dout0(n1861)
  );


  SyncRegister
  reg_C369
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1843),
    .dout0(n1848)
  );


  SyncRegister
  reg_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1272),
    .dout0(n1273)
  );


  SyncRegister
  reg_C370
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1861),
    .dout0(n1862)
  );


  SyncRegister
  reg_C371
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1862),
    .dout0(n1911)
  );


  SyncRegister
  reg_C372
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1852),
    .dout0(n1855)
  );


  SyncRegister
  reg_C373
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1866),
    .dout0(n1870)
  );


  SyncRegister
  reg_C374
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1874),
    .din0(n1910)
  );


  SyncRegister
  reg_C375
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1882),
    .din0(n1911)
  );


  SyncRegister
  reg_C376
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1888),
    .din0(n1910)
  );


  SyncRegister
  reg_C377
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1882),
    .dout0(n1883)
  );


  SyncRegister
  reg_C378
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1874),
    .dout0(n1875)
  );


  SyncRegister
  reg_C379
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1875),
    .dout0(n1876)
  );


  SyncRegister
  reg_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1290),
    .dout0(n1291)
  );


  SyncRegister
  reg_C380
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1883),
    .dout0(n1884)
  );


  SyncRegister
  reg_C381
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1876),
    .dout0(n1877)
  );


  SyncRegister
  reg_C382
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1884),
    .dout0(n1885)
  );


  SyncRegister
  reg_C383
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1877),
    .dout0(n1878)
  );


  SyncRegister
  reg_C384
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1878),
    .dout0(n1879)
  );


  SyncRegister
  reg_C385
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1896),
    .dout0(n1897)
  );


  SyncRegister
  reg_C386
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1896),
    .dout0(n1903)
  );


  SyncRegister
  reg_C387
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1879),
    .dout0(n1880)
  );


  SyncRegister
  reg_C388
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1897),
    .dout0(n1898)
  );


  SyncRegister
  reg_C389
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1880),
    .dout0(n1881)
  );


  SyncRegister
  reg_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1273),
    .dout0(n1278)
  );


  SyncRegister
  reg_C390
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1898),
    .dout0(n1899)
  );


  SyncRegister
  reg_C391
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1881),
    .dout0(n1886)
  );


  SyncRegister
  reg_C392
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1899),
    .dout0(n1900)
  );


  SyncRegister
  reg_C393
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1900),
    .dout0(n1949)
  );


  SyncRegister
  reg_C394
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1890),
    .dout0(n1893)
  );


  SyncRegister
  reg_C395
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1904),
    .dout0(n1908)
  );


  SyncRegister
  reg_C396
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1912),
    .din0(n1948)
  );


  SyncRegister
  reg_C397
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1920),
    .din0(n1949)
  );


  SyncRegister
  reg_C398
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1926),
    .din0(n1948)
  );


  SyncRegister
  reg_C399
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1920),
    .dout0(n1921)
  );


  SyncRegister
  reg_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1230),
    .dout0(n1231)
  );


  SyncRegister
  reg_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1291),
    .dout0(n1292)
  );


  SyncRegister
  reg_C400
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1912),
    .dout0(n1913)
  );


  SyncRegister
  reg_C401
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1913),
    .dout0(n1914)
  );


  SyncRegister
  reg_C402
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1921),
    .dout0(n1922)
  );


  SyncRegister
  reg_C403
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1914),
    .dout0(n1915)
  );


  SyncRegister
  reg_C404
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1922),
    .dout0(n1923)
  );


  SyncRegister
  reg_C405
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1915),
    .dout0(n1916)
  );


  SyncRegister
  reg_C406
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1916),
    .dout0(n1917)
  );


  SyncRegister
  reg_C407
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1934),
    .dout0(n1935)
  );


  SyncRegister
  reg_C408
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1934),
    .dout0(n1941)
  );


  SyncRegister
  reg_C409
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1917),
    .dout0(n1918)
  );


  SyncRegister
  reg_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1292),
    .dout0(n1341)
  );


  SyncRegister
  reg_C410
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1935),
    .dout0(n1936)
  );


  SyncRegister
  reg_C411
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1918),
    .dout0(n1919)
  );


  SyncRegister
  reg_C412
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1936),
    .dout0(n1937)
  );


  SyncRegister
  reg_C413
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1919),
    .dout0(n1924)
  );


  SyncRegister
  reg_C414
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1937),
    .dout0(n1938)
  );


  SyncRegister
  reg_C415
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1938),
    .dout0(n1987)
  );


  SyncRegister
  reg_C416
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1928),
    .dout0(n1931)
  );


  SyncRegister
  reg_C417
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1942),
    .dout0(n1946)
  );


  SyncRegister
  reg_C418
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1950),
    .din0(n1986)
  );


  SyncRegister
  reg_C419
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1958),
    .din0(n1987)
  );


  SyncRegister
  reg_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1282),
    .dout0(n1285)
  );


  SyncRegister
  reg_C420
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1964),
    .din0(n1986)
  );


  SyncRegister
  reg_C421
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1958),
    .dout0(n1959)
  );


  SyncRegister
  reg_C422
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1950),
    .dout0(n1951)
  );


  SyncRegister
  reg_C423
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1951),
    .dout0(n1952)
  );


  SyncRegister
  reg_C424
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1959),
    .dout0(n1960)
  );


  SyncRegister
  reg_C425
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1952),
    .dout0(n1953)
  );


  SyncRegister
  reg_C426
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1960),
    .dout0(n1961)
  );


  SyncRegister
  reg_C427
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1953),
    .dout0(n1954)
  );


  SyncRegister
  reg_C428
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1954),
    .dout0(n1955)
  );


  SyncRegister
  reg_C429
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1972),
    .dout0(n1973)
  );


  SyncRegister
  reg_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1296),
    .dout0(n1300)
  );


  SyncRegister
  reg_C430
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1972),
    .dout0(n1979)
  );


  SyncRegister
  reg_C431
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1955),
    .dout0(n1956)
  );


  SyncRegister
  reg_C432
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1973),
    .dout0(n1974)
  );


  SyncRegister
  reg_C433
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1956),
    .dout0(n1957)
  );


  SyncRegister
  reg_C434
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1974),
    .dout0(n1975)
  );


  SyncRegister
  reg_C435
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1957),
    .dout0(n1962)
  );


  SyncRegister
  reg_C436
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1975),
    .dout0(n1976)
  );


  SyncRegister
  reg_C437
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1976),
    .dout0(n2025)
  );


  SyncRegister
  reg_C438
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1966),
    .dout0(n1969)
  );


  SyncRegister
  reg_C439
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1980),
    .dout0(n1984)
  );


  SyncRegister
  reg_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1304),
    .din0(n1340)
  );


  SyncRegister
  reg_C440
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1988),
    .din0(n2024)
  );


  SyncRegister
  reg_C441
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1996),
    .din0(n2025)
  );


  SyncRegister
  reg_C442
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2002),
    .din0(n2024)
  );


  SyncRegister
  reg_C443
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1996),
    .dout0(n1997)
  );


  SyncRegister
  reg_C444
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1988),
    .dout0(n1989)
  );


  SyncRegister
  reg_C445
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1989),
    .dout0(n1990)
  );


  SyncRegister
  reg_C446
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1997),
    .dout0(n1998)
  );


  SyncRegister
  reg_C447
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1990),
    .dout0(n1991)
  );


  SyncRegister
  reg_C448
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1998),
    .dout0(n1999)
  );


  SyncRegister
  reg_C449
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1991),
    .dout0(n1992)
  );


  SyncRegister
  reg_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1312),
    .din0(n1341)
  );


  SyncRegister
  reg_C450
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1992),
    .dout0(n1993)
  );


  SyncRegister
  reg_C451
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2010),
    .dout0(n2011)
  );


  SyncRegister
  reg_C452
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2010),
    .dout0(n2017)
  );


  SyncRegister
  reg_C453
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1993),
    .dout0(n1994)
  );


  SyncRegister
  reg_C454
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2011),
    .dout0(n2012)
  );


  SyncRegister
  reg_C455
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1994),
    .dout0(n1995)
  );


  SyncRegister
  reg_C456
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2012),
    .dout0(n2013)
  );


  SyncRegister
  reg_C457
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1995),
    .dout0(n2000)
  );


  SyncRegister
  reg_C458
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2013),
    .dout0(n2014)
  );


  SyncRegister
  reg_C459
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2014),
    .dout0(n2063)
  );


  SyncRegister
  reg_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1318),
    .din0(n1340)
  );


  SyncRegister
  reg_C460
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2004),
    .dout0(n2007)
  );


  SyncRegister
  reg_C461
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2018),
    .dout0(n2022)
  );


  SyncRegister
  reg_C462
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2026),
    .din0(n2062)
  );


  SyncRegister
  reg_C463
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2034),
    .din0(n2063)
  );


  SyncRegister
  reg_C464
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2040),
    .din0(n2062)
  );


  SyncRegister
  reg_C465
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2034),
    .dout0(n2035)
  );


  SyncRegister
  reg_C466
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2026),
    .dout0(n2027)
  );


  SyncRegister
  reg_C467
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2027),
    .dout0(n2028)
  );


  SyncRegister
  reg_C468
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2035),
    .dout0(n2036)
  );


  SyncRegister
  reg_C469
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2028),
    .dout0(n2029)
  );


  SyncRegister
  reg_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1312),
    .dout0(n1313)
  );


  SyncRegister
  reg_C470
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2036),
    .dout0(n2037)
  );


  SyncRegister
  reg_C471
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2029),
    .dout0(n2030)
  );


  SyncRegister
  reg_C472
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2030),
    .dout0(n2031)
  );


  SyncRegister
  reg_C473
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2048),
    .dout0(n2049)
  );


  SyncRegister
  reg_C474
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2048),
    .dout0(n2055)
  );


  SyncRegister
  reg_C475
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2031),
    .dout0(n2032)
  );


  SyncRegister
  reg_C476
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2049),
    .dout0(n2050)
  );


  SyncRegister
  reg_C477
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2032),
    .dout0(n2033)
  );


  SyncRegister
  reg_C478
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2050),
    .dout0(n2051)
  );


  SyncRegister
  reg_C479
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2033),
    .dout0(n2038)
  );


  SyncRegister
  reg_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1304),
    .dout0(n1305)
  );


  SyncRegister
  reg_C480
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2051),
    .dout0(n2052)
  );


  SyncRegister
  reg_C481
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2052),
    .dout0(n2101)
  );


  SyncRegister
  reg_C482
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2042),
    .dout0(n2045)
  );


  SyncRegister
  reg_C483
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2056),
    .dout0(n2060)
  );


  SyncRegister
  reg_C484
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2064),
    .din0(n2100)
  );


  SyncRegister
  reg_C485
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2072),
    .din0(n2101)
  );


  SyncRegister
  reg_C486
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2078),
    .din0(n2100)
  );


  SyncRegister
  reg_C487
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2072),
    .dout0(n2073)
  );


  SyncRegister
  reg_C488
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2064),
    .dout0(n2065)
  );


  SyncRegister
  reg_C489
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2065),
    .dout0(n2066)
  );


  SyncRegister
  reg_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1305),
    .dout0(n1306)
  );


  SyncRegister
  reg_C490
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2073),
    .dout0(n2074)
  );


  SyncRegister
  reg_C491
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2066),
    .dout0(n2067)
  );


  SyncRegister
  reg_C492
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2074),
    .dout0(n2075)
  );


  SyncRegister
  reg_C493
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2067),
    .dout0(n2068)
  );


  SyncRegister
  reg_C494
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2068),
    .dout0(n2069)
  );


  SyncRegister
  reg_C495
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2086),
    .dout0(n2087)
  );


  SyncRegister
  reg_C496
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2086),
    .dout0(n2093)
  );


  SyncRegister
  reg_C497
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2069),
    .dout0(n2070)
  );


  SyncRegister
  reg_C498
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2087),
    .dout0(n2088)
  );


  SyncRegister
  reg_C499
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2070),
    .dout0(n2071)
  );


  SyncRegister
  reg_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1231),
    .dout0(n1232)
  );


  SyncRegister
  reg_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1313),
    .dout0(n1314)
  );


  SyncRegister
  reg_C500
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2088),
    .dout0(n2089)
  );


  SyncRegister
  reg_C501
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2071),
    .dout0(n2076)
  );


  SyncRegister
  reg_C502
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2089),
    .dout0(n2090)
  );


  SyncRegister
  reg_C503
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2090),
    .dout0(n2139)
  );


  SyncRegister
  reg_C504
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2080),
    .dout0(n2083)
  );


  SyncRegister
  reg_C505
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2094),
    .dout0(n2098)
  );


  SyncRegister
  reg_C506
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2102),
    .din0(n2138)
  );


  SyncRegister
  reg_C507
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2110),
    .din0(n2139)
  );


  SyncRegister
  reg_C508
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2116),
    .din0(n2138)
  );


  SyncRegister
  reg_C509
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2110),
    .dout0(n2111)
  );


  SyncRegister
  reg_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1306),
    .dout0(n1307)
  );


  SyncRegister
  reg_C510
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2102),
    .dout0(n2103)
  );


  SyncRegister
  reg_C511
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2103),
    .dout0(n2104)
  );


  SyncRegister
  reg_C512
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2111),
    .dout0(n2112)
  );


  SyncRegister
  reg_C513
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2104),
    .dout0(n2105)
  );


  SyncRegister
  reg_C514
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2112),
    .dout0(n2113)
  );


  SyncRegister
  reg_C515
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2105),
    .dout0(n2106)
  );


  SyncRegister
  reg_C516
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2106),
    .dout0(n2107)
  );


  SyncRegister
  reg_C517
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2124),
    .dout0(n2125)
  );


  SyncRegister
  reg_C518
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2124),
    .dout0(n2131)
  );


  SyncRegister
  reg_C519
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2107),
    .dout0(n2108)
  );


  SyncRegister
  reg_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1314),
    .dout0(n1315)
  );


  SyncRegister
  reg_C520
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2125),
    .dout0(n2126)
  );


  SyncRegister
  reg_C521
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2108),
    .dout0(n2109)
  );


  SyncRegister
  reg_C522
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2126),
    .dout0(n2127)
  );


  SyncRegister
  reg_C523
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2109),
    .dout0(n2114)
  );


  SyncRegister
  reg_C524
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2127),
    .dout0(n2128)
  );


  SyncRegister
  reg_C525
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2128),
    .dout0(n2177)
  );


  SyncRegister
  reg_C526
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2118),
    .dout0(n2121)
  );


  SyncRegister
  reg_C527
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2132),
    .dout0(n2136)
  );


  SyncRegister
  reg_C528
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2140),
    .din0(n2176)
  );


  SyncRegister
  reg_C529
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2148),
    .din0(n2177)
  );


  SyncRegister
  reg_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1307),
    .dout0(n1308)
  );


  SyncRegister
  reg_C530
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2154),
    .din0(n2176)
  );


  SyncRegister
  reg_C531
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2148),
    .dout0(n2149)
  );


  SyncRegister
  reg_C532
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2140),
    .dout0(n2141)
  );


  SyncRegister
  reg_C533
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2141),
    .dout0(n2142)
  );


  SyncRegister
  reg_C534
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2149),
    .dout0(n2150)
  );


  SyncRegister
  reg_C535
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2142),
    .dout0(n2143)
  );


  SyncRegister
  reg_C536
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2150),
    .dout0(n2151)
  );


  SyncRegister
  reg_C537
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2143),
    .dout0(n2144)
  );


  SyncRegister
  reg_C538
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2144),
    .dout0(n2145)
  );


  SyncRegister
  reg_C539
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2162),
    .dout0(n2163)
  );


  SyncRegister
  reg_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1308),
    .dout0(n1309)
  );


  SyncRegister
  reg_C540
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2162),
    .dout0(n2169)
  );


  SyncRegister
  reg_C541
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2145),
    .dout0(n2146)
  );


  SyncRegister
  reg_C542
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2163),
    .dout0(n2164)
  );


  SyncRegister
  reg_C543
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2146),
    .dout0(n2147)
  );


  SyncRegister
  reg_C544
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2164),
    .dout0(n2165)
  );


  SyncRegister
  reg_C545
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2147),
    .dout0(n2152)
  );


  SyncRegister
  reg_C546
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2165),
    .dout0(n2166)
  );


  SyncRegister
  reg_C547
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2166),
    .dout0(n2215)
  );


  SyncRegister
  reg_C548
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2156),
    .dout0(n2159)
  );


  SyncRegister
  reg_C549
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2170),
    .dout0(n2174)
  );


  SyncRegister
  reg_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1326),
    .dout0(n1327)
  );


  SyncRegister
  reg_C550
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2178),
    .din0(n2214)
  );


  SyncRegister
  reg_C551
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2186),
    .din0(n2215)
  );


  SyncRegister
  reg_C552
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2192),
    .din0(n2214)
  );


  SyncRegister
  reg_C553
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2186),
    .dout0(n2187)
  );


  SyncRegister
  reg_C554
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2178),
    .dout0(n2179)
  );


  SyncRegister
  reg_C555
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2179),
    .dout0(n2180)
  );


  SyncRegister
  reg_C556
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2187),
    .dout0(n2188)
  );


  SyncRegister
  reg_C557
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2180),
    .dout0(n2181)
  );


  SyncRegister
  reg_C558
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2188),
    .dout0(n2189)
  );


  SyncRegister
  reg_C559
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2181),
    .dout0(n2182)
  );


  SyncRegister
  reg_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1326),
    .dout0(n1333)
  );


  SyncRegister
  reg_C560
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2182),
    .dout0(n2183)
  );


  SyncRegister
  reg_C561
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2200),
    .dout0(n2201)
  );


  SyncRegister
  reg_C562
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2200),
    .dout0(n2207)
  );


  SyncRegister
  reg_C563
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2183),
    .dout0(n2184)
  );


  SyncRegister
  reg_C564
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2201),
    .dout0(n2202)
  );


  SyncRegister
  reg_C565
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2184),
    .dout0(n2185)
  );


  SyncRegister
  reg_C566
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2202),
    .dout0(n2203)
  );


  SyncRegister
  reg_C567
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2185),
    .dout0(n2190)
  );


  SyncRegister
  reg_C568
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2203),
    .dout0(n2204)
  );


  SyncRegister
  reg_C569
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2204),
    .dout0(n2253)
  );


  SyncRegister
  reg_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1309),
    .dout0(n1310)
  );


  SyncRegister
  reg_C570
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2194),
    .dout0(n2197)
  );


  SyncRegister
  reg_C571
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2208),
    .dout0(n2212)
  );


  SyncRegister
  reg_C572
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2216),
    .din0(n2252)
  );


  SyncRegister
  reg_C573
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2224),
    .din0(n2253)
  );


  SyncRegister
  reg_C574
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2230),
    .din0(n2252)
  );


  SyncRegister
  reg_C575
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2224),
    .dout0(n2225)
  );


  SyncRegister
  reg_C576
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2216),
    .dout0(n2217)
  );


  SyncRegister
  reg_C577
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2217),
    .dout0(n2218)
  );


  SyncRegister
  reg_C578
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2225),
    .dout0(n2226)
  );


  SyncRegister
  reg_C579
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2218),
    .dout0(n2219)
  );


  SyncRegister
  reg_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1327),
    .dout0(n1328)
  );


  SyncRegister
  reg_C580
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2226),
    .dout0(n2227)
  );


  SyncRegister
  reg_C581
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2219),
    .dout0(n2220)
  );


  SyncRegister
  reg_C582
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2220),
    .dout0(n2221)
  );


  SyncRegister
  reg_C583
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2238),
    .dout0(n2239)
  );


  SyncRegister
  reg_C584
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2238),
    .dout0(n2245)
  );


  SyncRegister
  reg_C585
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2221),
    .dout0(n2222)
  );


  SyncRegister
  reg_C586
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2239),
    .dout0(n2240)
  );


  SyncRegister
  reg_C587
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2222),
    .dout0(n2223)
  );


  SyncRegister
  reg_C588
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2240),
    .dout0(n2241)
  );


  SyncRegister
  reg_C589
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2223),
    .dout0(n2228)
  );


  SyncRegister
  reg_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1310),
    .dout0(n1311)
  );


  SyncRegister
  reg_C590
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2241),
    .dout0(n2242)
  );


  SyncRegister
  reg_C591
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2242),
    .dout0(n2291)
  );


  SyncRegister
  reg_C592
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2232),
    .dout0(n2235)
  );


  SyncRegister
  reg_C593
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2246),
    .dout0(n2250)
  );


  SyncRegister
  reg_C594
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2254),
    .din0(n2290)
  );


  SyncRegister
  reg_C595
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2262),
    .din0(n2291)
  );


  SyncRegister
  reg_C596
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2268),
    .din0(n2290)
  );


  SyncRegister
  reg_C597
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2262),
    .dout0(n2263)
  );


  SyncRegister
  reg_C598
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2254),
    .dout0(n2255)
  );


  SyncRegister
  reg_C599
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2255),
    .dout0(n2256)
  );


  SyncRegister
  reg_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1239),
    .dout0(n1240)
  );


  SyncRegister
  reg_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1328),
    .dout0(n1329)
  );


  SyncRegister
  reg_C600
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2263),
    .dout0(n2264)
  );


  SyncRegister
  reg_C601
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2256),
    .dout0(n2257)
  );


  SyncRegister
  reg_C602
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2264),
    .dout0(n2265)
  );


  SyncRegister
  reg_C603
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2257),
    .dout0(n2258)
  );


  SyncRegister
  reg_C604
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2258),
    .dout0(n2259)
  );


  SyncRegister
  reg_C605
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2276),
    .dout0(n2277)
  );


  SyncRegister
  reg_C606
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2276),
    .dout0(n2283)
  );


  SyncRegister
  reg_C607
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2259),
    .dout0(n2260)
  );


  SyncRegister
  reg_C608
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2277),
    .dout0(n2278)
  );


  SyncRegister
  reg_C609
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2260),
    .dout0(n2261)
  );


  SyncRegister
  reg_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1311),
    .dout0(n1316)
  );


  SyncRegister
  reg_C610
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2278),
    .dout0(n2279)
  );


  SyncRegister
  reg_C611
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2261),
    .dout0(n2266)
  );


  SyncRegister
  reg_C612
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2279),
    .dout0(n2280)
  );


  SyncRegister
  reg_C613
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2280),
    .dout0(n2329)
  );


  SyncRegister
  reg_C614
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2270),
    .dout0(n2273)
  );


  SyncRegister
  reg_C615
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2284),
    .dout0(n2288)
  );


  SyncRegister
  reg_C616
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2292),
    .din0(n2328)
  );


  SyncRegister
  reg_C617
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2300),
    .din0(n2329)
  );


  SyncRegister
  reg_C618
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2306),
    .din0(n2328)
  );


  SyncRegister
  reg_C619
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2300),
    .dout0(n2301)
  );


  SyncRegister
  reg_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1329),
    .dout0(n1330)
  );


  SyncRegister
  reg_C620
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2292),
    .dout0(n2293)
  );


  SyncRegister
  reg_C621
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2293),
    .dout0(n2294)
  );


  SyncRegister
  reg_C622
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2301),
    .dout0(n2302)
  );


  SyncRegister
  reg_C623
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2294),
    .dout0(n2295)
  );


  SyncRegister
  reg_C624
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2302),
    .dout0(n2303)
  );


  SyncRegister
  reg_C625
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2295),
    .dout0(n2296)
  );


  SyncRegister
  reg_C626
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2296),
    .dout0(n2297)
  );


  SyncRegister
  reg_C627
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2314),
    .dout0(n2315)
  );


  SyncRegister
  reg_C628
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2314),
    .dout0(n2321)
  );


  SyncRegister
  reg_C629
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2297),
    .dout0(n2298)
  );


  SyncRegister
  reg_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1330),
    .dout0(n1379)
  );


  SyncRegister
  reg_C630
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2315),
    .dout0(n2316)
  );


  SyncRegister
  reg_C631
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2298),
    .dout0(n2299)
  );


  SyncRegister
  reg_C632
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2316),
    .dout0(n2317)
  );


  SyncRegister
  reg_C633
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2299),
    .dout0(n2304)
  );


  SyncRegister
  reg_C634
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2317),
    .dout0(n2318)
  );


  SyncRegister
  reg_C635
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2318),
    .dout0(n2367)
  );


  SyncRegister
  reg_C636
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2308),
    .dout0(n2311)
  );


  SyncRegister
  reg_C637
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2322),
    .dout0(n2326)
  );


  SyncRegister
  reg_C638
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2330),
    .din0(n2366)
  );


  SyncRegister
  reg_C639
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2338),
    .din0(n2367)
  );


  SyncRegister
  reg_C64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1320),
    .dout0(n1323)
  );


  SyncRegister
  reg_C640
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2344),
    .din0(n2366)
  );


  SyncRegister
  reg_C641
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2338),
    .dout0(n2339)
  );


  SyncRegister
  reg_C642
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2330),
    .dout0(n2331)
  );


  SyncRegister
  reg_C643
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2331),
    .dout0(n2332)
  );


  SyncRegister
  reg_C644
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2339),
    .dout0(n2340)
  );


  SyncRegister
  reg_C645
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2332),
    .dout0(n2333)
  );


  SyncRegister
  reg_C646
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2340),
    .dout0(n2341)
  );


  SyncRegister
  reg_C647
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2333),
    .dout0(n2334)
  );


  SyncRegister
  reg_C648
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2334),
    .dout0(n2335)
  );


  SyncRegister
  reg_C649
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2352),
    .dout0(n2353)
  );


  SyncRegister
  reg_C65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1334),
    .dout0(n1338)
  );


  SyncRegister
  reg_C650
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2352),
    .dout0(n2359)
  );


  SyncRegister
  reg_C651
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2335),
    .dout0(n2336)
  );


  SyncRegister
  reg_C652
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2353),
    .dout0(n2354)
  );


  SyncRegister
  reg_C653
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2336),
    .dout0(n2337)
  );


  SyncRegister
  reg_C654
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2354),
    .dout0(n2355)
  );


  SyncRegister
  reg_C655
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2337),
    .dout0(n2342)
  );


  SyncRegister
  reg_C656
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2355),
    .dout0(n2356)
  );


  SyncRegister
  reg_C657
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2356),
    .dout0(n2405)
  );


  SyncRegister
  reg_C658
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2346),
    .dout0(n2349)
  );


  SyncRegister
  reg_C659
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2360),
    .dout0(n2364)
  );


  SyncRegister
  reg_C66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1342),
    .din0(n1378)
  );


  SyncRegister
  reg_C660
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2368),
    .din0(n2404)
  );


  SyncRegister
  reg_C661
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2376),
    .din0(n2405)
  );


  SyncRegister
  reg_C662
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2382),
    .din0(n2404)
  );


  SyncRegister
  reg_C663
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2376),
    .dout0(n2377)
  );


  SyncRegister
  reg_C664
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2368),
    .dout0(n2369)
  );


  SyncRegister
  reg_C665
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2369),
    .dout0(n2370)
  );


  SyncRegister
  reg_C666
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2377),
    .dout0(n2378)
  );


  SyncRegister
  reg_C667
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2370),
    .dout0(n2371)
  );


  SyncRegister
  reg_C668
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2378),
    .dout0(n2379)
  );


  SyncRegister
  reg_C669
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2371),
    .dout0(n2372)
  );


  SyncRegister
  reg_C67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1350),
    .din0(n1379)
  );


  SyncRegister
  reg_C670
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2372),
    .dout0(n2373)
  );


  SyncRegister
  reg_C671
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2390),
    .dout0(n2391)
  );


  SyncRegister
  reg_C672
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2390),
    .dout0(n2397)
  );


  SyncRegister
  reg_C673
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2373),
    .dout0(n2374)
  );


  SyncRegister
  reg_C674
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2391),
    .dout0(n2392)
  );


  SyncRegister
  reg_C675
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2374),
    .dout0(n2375)
  );


  SyncRegister
  reg_C676
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2392),
    .dout0(n2393)
  );


  SyncRegister
  reg_C677
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2375),
    .dout0(n2380)
  );


  SyncRegister
  reg_C678
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2393),
    .dout0(n2394)
  );


  SyncRegister
  reg_C679
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2394),
    .dout0(n2443)
  );


  SyncRegister
  reg_C68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1356),
    .din0(n1378)
  );


  SyncRegister
  reg_C680
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2384),
    .dout0(n2387)
  );


  SyncRegister
  reg_C681
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2398),
    .dout0(n2402)
  );


  SyncRegister
  reg_C682
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2406),
    .din0(n2442)
  );


  SyncRegister
  reg_C683
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2414),
    .din0(n2443)
  );


  SyncRegister
  reg_C684
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2420),
    .din0(n2442)
  );


  SyncRegister
  reg_C685
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2414),
    .dout0(n2415)
  );


  SyncRegister
  reg_C686
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2406),
    .dout0(n2407)
  );


  SyncRegister
  reg_C687
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2407),
    .dout0(n2408)
  );


  SyncRegister
  reg_C688
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2415),
    .dout0(n2416)
  );


  SyncRegister
  reg_C689
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2408),
    .dout0(n2409)
  );


  SyncRegister
  reg_C69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1350),
    .dout0(n1351)
  );


  SyncRegister
  reg_C690
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2416),
    .dout0(n2417)
  );


  SyncRegister
  reg_C691
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2409),
    .dout0(n2410)
  );


  SyncRegister
  reg_C692
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2410),
    .dout0(n2411)
  );


  SyncRegister
  reg_C693
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2428),
    .dout0(n2429)
  );


  SyncRegister
  reg_C694
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2428),
    .dout0(n2435)
  );


  SyncRegister
  reg_C695
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2411),
    .dout0(n2412)
  );


  SyncRegister
  reg_C696
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2429),
    .dout0(n2430)
  );


  SyncRegister
  reg_C697
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2412),
    .dout0(n2413)
  );


  SyncRegister
  reg_C698
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2430),
    .dout0(n2431)
  );


  SyncRegister
  reg_C699
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2413),
    .dout0(n2418)
  );


  SyncRegister
  reg_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1232),
    .dout0(n1233)
  );


  SyncRegister
  reg_C70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1342),
    .dout0(n1343)
  );


  SyncRegister
  reg_C700
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2431),
    .dout0(n2432)
  );


  SyncRegister
  reg_C701
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2432),
    .dout0(n2449)
  );


  SyncRegister
  reg_C702
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2422),
    .dout0(n2425)
  );


  SyncRegister
  reg_C703
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2436),
    .dout0(n2440)
  );


  SyncRegister
  reg_C71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1343),
    .dout0(n1344)
  );


  SyncRegister
  reg_C72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1351),
    .dout0(n1352)
  );


  SyncRegister
  reg_C73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1344),
    .dout0(n1345)
  );


  SyncRegister
  reg_C74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1352),
    .dout0(n1353)
  );


  SyncRegister
  reg_C75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1345),
    .dout0(n1346)
  );


  SyncRegister
  reg_C76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1346),
    .dout0(n1347)
  );


  SyncRegister
  reg_C77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1364),
    .dout0(n1365)
  );


  SyncRegister
  reg_C78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1364),
    .dout0(n1371)
  );


  SyncRegister
  reg_C79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1347),
    .dout0(n1348)
  );


  SyncRegister
  reg_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1240),
    .dout0(n1241)
  );


  SyncRegister
  reg_C80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1365),
    .dout0(n1366)
  );


  SyncRegister
  reg_C81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1348),
    .dout0(n1349)
  );


  SyncRegister
  reg_C82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1366),
    .dout0(n1367)
  );


  SyncRegister
  reg_C83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1349),
    .dout0(n1354)
  );


  SyncRegister
  reg_C84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1367),
    .dout0(n1368)
  );


  SyncRegister
  reg_C85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1368),
    .dout0(n1417)
  );


  SyncRegister
  reg_C86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1358),
    .dout0(n1361)
  );


  SyncRegister
  reg_C87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1372),
    .dout0(n1376)
  );


  SyncRegister
  reg_C88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1380),
    .din0(n1416)
  );


  SyncRegister
  reg_C89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1388),
    .din0(n1417)
  );


  SyncRegister
  reg_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1233),
    .dout0(n1234)
  );


  SyncRegister
  reg_C90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1394),
    .din0(n1416)
  );


  SyncRegister
  reg_C91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1388),
    .dout0(n1389)
  );


  SyncRegister
  reg_C92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1380),
    .dout0(n1381)
  );


  SyncRegister
  reg_C93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1381),
    .dout0(n1382)
  );


  SyncRegister
  reg_C94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1389),
    .dout0(n1390)
  );


  SyncRegister
  reg_C95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1382),
    .dout0(n1383)
  );


  SyncRegister
  reg_C96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1390),
    .dout0(n1391)
  );


  SyncRegister
  reg_C97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1383),
    .dout0(n1384)
  );


  SyncRegister
  reg_C98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1384),
    .dout0(n1385)
  );


  SyncRegister
  reg_C99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1402),
    .dout0(n1403)
  );


  SyncRegister
  reg_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n0),
    .din0(n2444)
  );


  SyncRegister
  reg_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2445),
    .dout0(n8)
  );


  SyncRegister
  reg_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n4),
    .dout0(n5)
  );


  SyncRegister
  reg_D100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n172),
    .dout0(n179)
  );


  SyncRegister
  reg_D101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n155),
    .dout0(n156)
  );


  SyncRegister
  reg_D102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n173),
    .dout0(n174)
  );


  SyncRegister
  reg_D103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n156),
    .dout0(n157)
  );


  SyncRegister
  reg_D104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n174),
    .dout0(n175)
  );


  SyncRegister
  reg_D105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n157),
    .dout0(n162)
  );


  SyncRegister
  reg_D106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n175),
    .dout0(n176)
  );


  SyncRegister
  reg_D107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n176),
    .dout0(n225)
  );


  SyncRegister
  reg_D108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n166),
    .dout0(n169)
  );


  SyncRegister
  reg_D109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n180),
    .dout0(n184)
  );


  SyncRegister
  reg_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n22),
    .dout0(n23)
  );


  SyncRegister
  reg_D110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n188),
    .din0(n224)
  );


  SyncRegister
  reg_D111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n196),
    .din0(n225)
  );


  SyncRegister
  reg_D112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n202),
    .din0(n224)
  );


  SyncRegister
  reg_D113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n196),
    .dout0(n197)
  );


  SyncRegister
  reg_D114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n188),
    .dout0(n189)
  );


  SyncRegister
  reg_D115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n189),
    .dout0(n190)
  );


  SyncRegister
  reg_D116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n197),
    .dout0(n198)
  );


  SyncRegister
  reg_D117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n190),
    .dout0(n191)
  );


  SyncRegister
  reg_D118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n198),
    .dout0(n199)
  );


  SyncRegister
  reg_D119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n191),
    .dout0(n192)
  );


  SyncRegister
  reg_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n22),
    .dout0(n29)
  );


  SyncRegister
  reg_D120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n192),
    .dout0(n193)
  );


  SyncRegister
  reg_D121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n210),
    .dout0(n211)
  );


  SyncRegister
  reg_D122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n210),
    .dout0(n217)
  );


  SyncRegister
  reg_D123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n193),
    .dout0(n194)
  );


  SyncRegister
  reg_D124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n211),
    .dout0(n212)
  );


  SyncRegister
  reg_D125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n194),
    .dout0(n195)
  );


  SyncRegister
  reg_D126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n212),
    .dout0(n213)
  );


  SyncRegister
  reg_D127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n195),
    .dout0(n200)
  );


  SyncRegister
  reg_D128
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n213),
    .dout0(n214)
  );


  SyncRegister
  reg_D129
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n214),
    .dout0(n263)
  );


  SyncRegister
  reg_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n5),
    .dout0(n6)
  );


  SyncRegister
  reg_D130
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n204),
    .dout0(n207)
  );


  SyncRegister
  reg_D131
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n218),
    .dout0(n222)
  );


  SyncRegister
  reg_D132
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n226),
    .din0(n262)
  );


  SyncRegister
  reg_D133
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n234),
    .din0(n263)
  );


  SyncRegister
  reg_D134
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n240),
    .din0(n262)
  );


  SyncRegister
  reg_D135
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n234),
    .dout0(n235)
  );


  SyncRegister
  reg_D136
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n226),
    .dout0(n227)
  );


  SyncRegister
  reg_D137
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n227),
    .dout0(n228)
  );


  SyncRegister
  reg_D138
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n235),
    .dout0(n236)
  );


  SyncRegister
  reg_D139
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n228),
    .dout0(n229)
  );


  SyncRegister
  reg_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n23),
    .dout0(n24)
  );


  SyncRegister
  reg_D140
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n236),
    .dout0(n237)
  );


  SyncRegister
  reg_D141
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n229),
    .dout0(n230)
  );


  SyncRegister
  reg_D142
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n230),
    .dout0(n231)
  );


  SyncRegister
  reg_D143
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n248),
    .dout0(n249)
  );


  SyncRegister
  reg_D144
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n248),
    .dout0(n255)
  );


  SyncRegister
  reg_D145
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n231),
    .dout0(n232)
  );


  SyncRegister
  reg_D146
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n249),
    .dout0(n250)
  );


  SyncRegister
  reg_D147
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n232),
    .dout0(n233)
  );


  SyncRegister
  reg_D148
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n250),
    .dout0(n251)
  );


  SyncRegister
  reg_D149
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n233),
    .dout0(n238)
  );


  SyncRegister
  reg_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n6),
    .dout0(n7)
  );


  SyncRegister
  reg_D150
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n251),
    .dout0(n252)
  );


  SyncRegister
  reg_D151
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n252),
    .dout0(n301)
  );


  SyncRegister
  reg_D152
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n242),
    .dout0(n245)
  );


  SyncRegister
  reg_D153
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n256),
    .dout0(n260)
  );


  SyncRegister
  reg_D154
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n264),
    .din0(n300)
  );


  SyncRegister
  reg_D155
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n272),
    .din0(n301)
  );


  SyncRegister
  reg_D156
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n278),
    .din0(n300)
  );


  SyncRegister
  reg_D157
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n272),
    .dout0(n273)
  );


  SyncRegister
  reg_D158
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n264),
    .dout0(n265)
  );


  SyncRegister
  reg_D159
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n265),
    .dout0(n266)
  );


  SyncRegister
  reg_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n24),
    .dout0(n25)
  );


  SyncRegister
  reg_D160
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n273),
    .dout0(n274)
  );


  SyncRegister
  reg_D161
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n266),
    .dout0(n267)
  );


  SyncRegister
  reg_D162
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n274),
    .dout0(n275)
  );


  SyncRegister
  reg_D163
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n267),
    .dout0(n268)
  );


  SyncRegister
  reg_D164
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n268),
    .dout0(n269)
  );


  SyncRegister
  reg_D165
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n286),
    .dout0(n287)
  );


  SyncRegister
  reg_D166
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n286),
    .dout0(n293)
  );


  SyncRegister
  reg_D167
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n269),
    .dout0(n270)
  );


  SyncRegister
  reg_D168
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n287),
    .dout0(n288)
  );


  SyncRegister
  reg_D169
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n270),
    .dout0(n271)
  );


  SyncRegister
  reg_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n12),
    .din0(n7)
  );


  SyncRegister
  reg_D170
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n288),
    .dout0(n289)
  );


  SyncRegister
  reg_D171
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n271),
    .dout0(n276)
  );


  SyncRegister
  reg_D172
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n289),
    .dout0(n290)
  );


  SyncRegister
  reg_D173
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n290),
    .dout0(n339)
  );


  SyncRegister
  reg_D174
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n280),
    .dout0(n283)
  );


  SyncRegister
  reg_D175
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n294),
    .dout0(n298)
  );


  SyncRegister
  reg_D176
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n302),
    .din0(n338)
  );


  SyncRegister
  reg_D177
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n310),
    .din0(n339)
  );


  SyncRegister
  reg_D178
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n316),
    .din0(n338)
  );


  SyncRegister
  reg_D179
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n310),
    .dout0(n311)
  );


  SyncRegister
  reg_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n25),
    .dout0(n26)
  );


  SyncRegister
  reg_D180
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n302),
    .dout0(n303)
  );


  SyncRegister
  reg_D181
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n303),
    .dout0(n304)
  );


  SyncRegister
  reg_D182
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n311),
    .dout0(n312)
  );


  SyncRegister
  reg_D183
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n304),
    .dout0(n305)
  );


  SyncRegister
  reg_D184
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n312),
    .dout0(n313)
  );


  SyncRegister
  reg_D185
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n305),
    .dout0(n306)
  );


  SyncRegister
  reg_D186
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n306),
    .dout0(n307)
  );


  SyncRegister
  reg_D187
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n324),
    .dout0(n325)
  );


  SyncRegister
  reg_D188
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n324),
    .dout0(n331)
  );


  SyncRegister
  reg_D189
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n307),
    .dout0(n308)
  );


  SyncRegister
  reg_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n26),
    .dout0(n73)
  );


  SyncRegister
  reg_D190
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n325),
    .dout0(n326)
  );


  SyncRegister
  reg_D191
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n308),
    .dout0(n309)
  );


  SyncRegister
  reg_D192
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n326),
    .dout0(n327)
  );


  SyncRegister
  reg_D193
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n309),
    .dout0(n314)
  );


  SyncRegister
  reg_D194
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n327),
    .dout0(n328)
  );


  SyncRegister
  reg_D195
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n328),
    .dout0(n377)
  );


  SyncRegister
  reg_D196
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n318),
    .dout0(n321)
  );


  SyncRegister
  reg_D197
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n332),
    .dout0(n336)
  );


  SyncRegister
  reg_D198
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n340),
    .din0(n376)
  );


  SyncRegister
  reg_D199
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n348),
    .din0(n377)
  );


  SyncRegister
  reg_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n14),
    .din0(n2444)
  );


  SyncRegister
  reg_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n16),
    .dout0(n19)
  );


  SyncRegister
  reg_D200
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n354),
    .din0(n376)
  );


  SyncRegister
  reg_D201
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n348),
    .dout0(n349)
  );


  SyncRegister
  reg_D202
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n340),
    .dout0(n341)
  );


  SyncRegister
  reg_D203
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n341),
    .dout0(n342)
  );


  SyncRegister
  reg_D204
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n349),
    .dout0(n350)
  );


  SyncRegister
  reg_D205
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n342),
    .dout0(n343)
  );


  SyncRegister
  reg_D206
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n350),
    .dout0(n351)
  );


  SyncRegister
  reg_D207
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n343),
    .dout0(n344)
  );


  SyncRegister
  reg_D208
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n344),
    .dout0(n345)
  );


  SyncRegister
  reg_D209
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n362),
    .dout0(n363)
  );


  SyncRegister
  reg_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n30),
    .dout0(n34)
  );


  SyncRegister
  reg_D210
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n362),
    .dout0(n369)
  );


  SyncRegister
  reg_D211
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n345),
    .dout0(n346)
  );


  SyncRegister
  reg_D212
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n363),
    .dout0(n364)
  );


  SyncRegister
  reg_D213
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n346),
    .dout0(n347)
  );


  SyncRegister
  reg_D214
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n364),
    .dout0(n365)
  );


  SyncRegister
  reg_D215
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n347),
    .dout0(n352)
  );


  SyncRegister
  reg_D216
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n365),
    .dout0(n366)
  );


  SyncRegister
  reg_D217
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n366),
    .dout0(n415)
  );


  SyncRegister
  reg_D218
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n356),
    .dout0(n359)
  );


  SyncRegister
  reg_D219
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n370),
    .dout0(n374)
  );


  SyncRegister
  reg_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n36),
    .din0(n72)
  );


  SyncRegister
  reg_D220
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n378),
    .din0(n414)
  );


  SyncRegister
  reg_D221
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n386),
    .din0(n415)
  );


  SyncRegister
  reg_D222
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n392),
    .din0(n414)
  );


  SyncRegister
  reg_D223
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n386),
    .dout0(n387)
  );


  SyncRegister
  reg_D224
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n378),
    .dout0(n379)
  );


  SyncRegister
  reg_D225
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n379),
    .dout0(n380)
  );


  SyncRegister
  reg_D226
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n387),
    .dout0(n388)
  );


  SyncRegister
  reg_D227
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n380),
    .dout0(n381)
  );


  SyncRegister
  reg_D228
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n388),
    .dout0(n389)
  );


  SyncRegister
  reg_D229
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n381),
    .dout0(n382)
  );


  SyncRegister
  reg_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n44),
    .din0(n73)
  );


  SyncRegister
  reg_D230
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n382),
    .dout0(n383)
  );


  SyncRegister
  reg_D231
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n400),
    .dout0(n401)
  );


  SyncRegister
  reg_D232
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n400),
    .dout0(n407)
  );


  SyncRegister
  reg_D233
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n383),
    .dout0(n384)
  );


  SyncRegister
  reg_D234
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n401),
    .dout0(n402)
  );


  SyncRegister
  reg_D235
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n384),
    .dout0(n385)
  );


  SyncRegister
  reg_D236
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n402),
    .dout0(n403)
  );


  SyncRegister
  reg_D237
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n385),
    .dout0(n390)
  );


  SyncRegister
  reg_D238
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n403),
    .dout0(n404)
  );


  SyncRegister
  reg_D239
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n404),
    .dout0(n453)
  );


  SyncRegister
  reg_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n50),
    .din0(n72)
  );


  SyncRegister
  reg_D240
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n394),
    .dout0(n397)
  );


  SyncRegister
  reg_D241
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n408),
    .dout0(n412)
  );


  SyncRegister
  reg_D242
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n416),
    .din0(n452)
  );


  SyncRegister
  reg_D243
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n424),
    .din0(n453)
  );


  SyncRegister
  reg_D244
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n430),
    .din0(n452)
  );


  SyncRegister
  reg_D245
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n424),
    .dout0(n425)
  );


  SyncRegister
  reg_D246
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n416),
    .dout0(n417)
  );


  SyncRegister
  reg_D247
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n417),
    .dout0(n418)
  );


  SyncRegister
  reg_D248
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n425),
    .dout0(n426)
  );


  SyncRegister
  reg_D249
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n418),
    .dout0(n419)
  );


  SyncRegister
  reg_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n44),
    .dout0(n45)
  );


  SyncRegister
  reg_D250
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n426),
    .dout0(n427)
  );


  SyncRegister
  reg_D251
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n419),
    .dout0(n420)
  );


  SyncRegister
  reg_D252
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n420),
    .dout0(n421)
  );


  SyncRegister
  reg_D253
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n438),
    .dout0(n439)
  );


  SyncRegister
  reg_D254
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n438),
    .dout0(n445)
  );


  SyncRegister
  reg_D255
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n421),
    .dout0(n422)
  );


  SyncRegister
  reg_D256
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n439),
    .dout0(n440)
  );


  SyncRegister
  reg_D257
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n422),
    .dout0(n423)
  );


  SyncRegister
  reg_D258
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n440),
    .dout0(n441)
  );


  SyncRegister
  reg_D259
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n423),
    .dout0(n428)
  );


  SyncRegister
  reg_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n36),
    .dout0(n37)
  );


  SyncRegister
  reg_D260
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n441),
    .dout0(n442)
  );


  SyncRegister
  reg_D261
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n442),
    .dout0(n491)
  );


  SyncRegister
  reg_D262
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n432),
    .dout0(n435)
  );


  SyncRegister
  reg_D263
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n446),
    .dout0(n450)
  );


  SyncRegister
  reg_D264
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n454),
    .din0(n490)
  );


  SyncRegister
  reg_D265
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n462),
    .din0(n491)
  );


  SyncRegister
  reg_D266
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n468),
    .din0(n490)
  );


  SyncRegister
  reg_D267
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n462),
    .dout0(n463)
  );


  SyncRegister
  reg_D268
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n454),
    .dout0(n455)
  );


  SyncRegister
  reg_D269
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n455),
    .dout0(n456)
  );


  SyncRegister
  reg_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n37),
    .dout0(n38)
  );


  SyncRegister
  reg_D270
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n463),
    .dout0(n464)
  );


  SyncRegister
  reg_D271
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n456),
    .dout0(n457)
  );


  SyncRegister
  reg_D272
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n464),
    .dout0(n465)
  );


  SyncRegister
  reg_D273
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n457),
    .dout0(n458)
  );


  SyncRegister
  reg_D274
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n458),
    .dout0(n459)
  );


  SyncRegister
  reg_D275
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n476),
    .dout0(n477)
  );


  SyncRegister
  reg_D276
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n476),
    .dout0(n483)
  );


  SyncRegister
  reg_D277
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n459),
    .dout0(n460)
  );


  SyncRegister
  reg_D278
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n477),
    .dout0(n478)
  );


  SyncRegister
  reg_D279
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n460),
    .dout0(n461)
  );


  SyncRegister
  reg_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n45),
    .dout0(n46)
  );


  SyncRegister
  reg_D280
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n478),
    .dout0(n479)
  );


  SyncRegister
  reg_D281
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n461),
    .dout0(n466)
  );


  SyncRegister
  reg_D282
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n479),
    .dout0(n480)
  );


  SyncRegister
  reg_D283
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n480),
    .dout0(n529)
  );


  SyncRegister
  reg_D284
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n470),
    .dout0(n473)
  );


  SyncRegister
  reg_D285
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n484),
    .dout0(n488)
  );


  SyncRegister
  reg_D286
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n492),
    .din0(n528)
  );


  SyncRegister
  reg_D287
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n500),
    .din0(n529)
  );


  SyncRegister
  reg_D288
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n506),
    .din0(n528)
  );


  SyncRegister
  reg_D289
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n500),
    .dout0(n501)
  );


  SyncRegister
  reg_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n38),
    .dout0(n39)
  );


  SyncRegister
  reg_D290
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n492),
    .dout0(n493)
  );


  SyncRegister
  reg_D291
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n493),
    .dout0(n494)
  );


  SyncRegister
  reg_D292
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n501),
    .dout0(n502)
  );


  SyncRegister
  reg_D293
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n494),
    .dout0(n495)
  );


  SyncRegister
  reg_D294
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n502),
    .dout0(n503)
  );


  SyncRegister
  reg_D295
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n495),
    .dout0(n496)
  );


  SyncRegister
  reg_D296
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n496),
    .dout0(n497)
  );


  SyncRegister
  reg_D297
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n514),
    .dout0(n515)
  );


  SyncRegister
  reg_D298
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n514),
    .dout0(n521)
  );


  SyncRegister
  reg_D299
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n497),
    .dout0(n498)
  );


  SyncRegister
  reg_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n8),
    .dout0(n9)
  );


  SyncRegister
  reg_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n46),
    .dout0(n47)
  );


  SyncRegister
  reg_D300
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n515),
    .dout0(n516)
  );


  SyncRegister
  reg_D301
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n498),
    .dout0(n499)
  );


  SyncRegister
  reg_D302
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n516),
    .dout0(n517)
  );


  SyncRegister
  reg_D303
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n499),
    .dout0(n504)
  );


  SyncRegister
  reg_D304
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n517),
    .dout0(n518)
  );


  SyncRegister
  reg_D305
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n518),
    .dout0(n567)
  );


  SyncRegister
  reg_D306
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n508),
    .dout0(n511)
  );


  SyncRegister
  reg_D307
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n522),
    .dout0(n526)
  );


  SyncRegister
  reg_D308
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n530),
    .din0(n566)
  );


  SyncRegister
  reg_D309
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n538),
    .din0(n567)
  );


  SyncRegister
  reg_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n39),
    .dout0(n40)
  );


  SyncRegister
  reg_D310
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n544),
    .din0(n566)
  );


  SyncRegister
  reg_D311
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n538),
    .dout0(n539)
  );


  SyncRegister
  reg_D312
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n530),
    .dout0(n531)
  );


  SyncRegister
  reg_D313
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n531),
    .dout0(n532)
  );


  SyncRegister
  reg_D314
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n539),
    .dout0(n540)
  );


  SyncRegister
  reg_D315
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n532),
    .dout0(n533)
  );


  SyncRegister
  reg_D316
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n540),
    .dout0(n541)
  );


  SyncRegister
  reg_D317
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n533),
    .dout0(n534)
  );


  SyncRegister
  reg_D318
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n534),
    .dout0(n535)
  );


  SyncRegister
  reg_D319
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n552),
    .dout0(n553)
  );


  SyncRegister
  reg_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n40),
    .dout0(n41)
  );


  SyncRegister
  reg_D320
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n552),
    .dout0(n559)
  );


  SyncRegister
  reg_D321
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n535),
    .dout0(n536)
  );


  SyncRegister
  reg_D322
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n553),
    .dout0(n554)
  );


  SyncRegister
  reg_D323
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n536),
    .dout0(n537)
  );


  SyncRegister
  reg_D324
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n554),
    .dout0(n555)
  );


  SyncRegister
  reg_D325
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n537),
    .dout0(n542)
  );


  SyncRegister
  reg_D326
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n555),
    .dout0(n556)
  );


  SyncRegister
  reg_D327
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n556),
    .dout0(n605)
  );


  SyncRegister
  reg_D328
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n546),
    .dout0(n549)
  );


  SyncRegister
  reg_D329
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n560),
    .dout0(n564)
  );


  SyncRegister
  reg_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n58),
    .dout0(n59)
  );


  SyncRegister
  reg_D330
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n568),
    .din0(n604)
  );


  SyncRegister
  reg_D331
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n576),
    .din0(n605)
  );


  SyncRegister
  reg_D332
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n582),
    .din0(n604)
  );


  SyncRegister
  reg_D333
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n576),
    .dout0(n577)
  );


  SyncRegister
  reg_D334
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n568),
    .dout0(n569)
  );


  SyncRegister
  reg_D335
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n569),
    .dout0(n570)
  );


  SyncRegister
  reg_D336
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n577),
    .dout0(n578)
  );


  SyncRegister
  reg_D337
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n570),
    .dout0(n571)
  );


  SyncRegister
  reg_D338
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n578),
    .dout0(n579)
  );


  SyncRegister
  reg_D339
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n571),
    .dout0(n572)
  );


  SyncRegister
  reg_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n58),
    .dout0(n65)
  );


  SyncRegister
  reg_D340
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n572),
    .dout0(n573)
  );


  SyncRegister
  reg_D341
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n590),
    .dout0(n591)
  );


  SyncRegister
  reg_D342
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n590),
    .dout0(n597)
  );


  SyncRegister
  reg_D343
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n573),
    .dout0(n574)
  );


  SyncRegister
  reg_D344
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n591),
    .dout0(n592)
  );


  SyncRegister
  reg_D345
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n574),
    .dout0(n575)
  );


  SyncRegister
  reg_D346
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n592),
    .dout0(n593)
  );


  SyncRegister
  reg_D347
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n575),
    .dout0(n580)
  );


  SyncRegister
  reg_D348
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n593),
    .dout0(n594)
  );


  SyncRegister
  reg_D349
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n594),
    .dout0(n643)
  );


  SyncRegister
  reg_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n41),
    .dout0(n42)
  );


  SyncRegister
  reg_D350
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n584),
    .dout0(n587)
  );


  SyncRegister
  reg_D351
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n598),
    .dout0(n602)
  );


  SyncRegister
  reg_D352
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n606),
    .din0(n642)
  );


  SyncRegister
  reg_D353
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n614),
    .din0(n643)
  );


  SyncRegister
  reg_D354
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n620),
    .din0(n642)
  );


  SyncRegister
  reg_D355
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n614),
    .dout0(n615)
  );


  SyncRegister
  reg_D356
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n606),
    .dout0(n607)
  );


  SyncRegister
  reg_D357
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n607),
    .dout0(n608)
  );


  SyncRegister
  reg_D358
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n615),
    .dout0(n616)
  );


  SyncRegister
  reg_D359
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n608),
    .dout0(n609)
  );


  SyncRegister
  reg_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n59),
    .dout0(n60)
  );


  SyncRegister
  reg_D360
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n616),
    .dout0(n617)
  );


  SyncRegister
  reg_D361
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n609),
    .dout0(n610)
  );


  SyncRegister
  reg_D362
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n610),
    .dout0(n611)
  );


  SyncRegister
  reg_D363
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n628),
    .dout0(n629)
  );


  SyncRegister
  reg_D364
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n628),
    .dout0(n635)
  );


  SyncRegister
  reg_D365
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n611),
    .dout0(n612)
  );


  SyncRegister
  reg_D366
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n629),
    .dout0(n630)
  );


  SyncRegister
  reg_D367
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n612),
    .dout0(n613)
  );


  SyncRegister
  reg_D368
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n630),
    .dout0(n631)
  );


  SyncRegister
  reg_D369
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n613),
    .dout0(n618)
  );


  SyncRegister
  reg_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n42),
    .dout0(n43)
  );


  SyncRegister
  reg_D370
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n631),
    .dout0(n632)
  );


  SyncRegister
  reg_D371
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n632),
    .dout0(n681)
  );


  SyncRegister
  reg_D372
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n622),
    .dout0(n625)
  );


  SyncRegister
  reg_D373
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n636),
    .dout0(n640)
  );


  SyncRegister
  reg_D374
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n644),
    .din0(n680)
  );


  SyncRegister
  reg_D375
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n652),
    .din0(n681)
  );


  SyncRegister
  reg_D376
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n658),
    .din0(n680)
  );


  SyncRegister
  reg_D377
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n652),
    .dout0(n653)
  );


  SyncRegister
  reg_D378
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n644),
    .dout0(n645)
  );


  SyncRegister
  reg_D379
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n645),
    .dout0(n646)
  );


  SyncRegister
  reg_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n60),
    .dout0(n61)
  );


  SyncRegister
  reg_D380
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n653),
    .dout0(n654)
  );


  SyncRegister
  reg_D381
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n646),
    .dout0(n647)
  );


  SyncRegister
  reg_D382
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n654),
    .dout0(n655)
  );


  SyncRegister
  reg_D383
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n647),
    .dout0(n648)
  );


  SyncRegister
  reg_D384
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n648),
    .dout0(n649)
  );


  SyncRegister
  reg_D385
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n666),
    .dout0(n667)
  );


  SyncRegister
  reg_D386
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n666),
    .dout0(n673)
  );


  SyncRegister
  reg_D387
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n649),
    .dout0(n650)
  );


  SyncRegister
  reg_D388
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n667),
    .dout0(n668)
  );


  SyncRegister
  reg_D389
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n650),
    .dout0(n651)
  );


  SyncRegister
  reg_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n43),
    .dout0(n48)
  );


  SyncRegister
  reg_D390
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n668),
    .dout0(n669)
  );


  SyncRegister
  reg_D391
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n651),
    .dout0(n656)
  );


  SyncRegister
  reg_D392
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n669),
    .dout0(n670)
  );


  SyncRegister
  reg_D393
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n670),
    .dout0(n719)
  );


  SyncRegister
  reg_D394
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n660),
    .dout0(n663)
  );


  SyncRegister
  reg_D395
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n674),
    .dout0(n678)
  );


  SyncRegister
  reg_D396
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n682),
    .din0(n718)
  );


  SyncRegister
  reg_D397
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n690),
    .din0(n719)
  );


  SyncRegister
  reg_D398
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n696),
    .din0(n718)
  );


  SyncRegister
  reg_D399
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n690),
    .dout0(n691)
  );


  SyncRegister
  reg_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n0),
    .dout0(n1)
  );


  SyncRegister
  reg_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n61),
    .dout0(n62)
  );


  SyncRegister
  reg_D400
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n682),
    .dout0(n683)
  );


  SyncRegister
  reg_D401
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n683),
    .dout0(n684)
  );


  SyncRegister
  reg_D402
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n691),
    .dout0(n692)
  );


  SyncRegister
  reg_D403
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n684),
    .dout0(n685)
  );


  SyncRegister
  reg_D404
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n692),
    .dout0(n693)
  );


  SyncRegister
  reg_D405
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n685),
    .dout0(n686)
  );


  SyncRegister
  reg_D406
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n686),
    .dout0(n687)
  );


  SyncRegister
  reg_D407
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n704),
    .dout0(n705)
  );


  SyncRegister
  reg_D408
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n704),
    .dout0(n711)
  );


  SyncRegister
  reg_D409
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n687),
    .dout0(n688)
  );


  SyncRegister
  reg_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n111),
    .din0(n62)
  );


  SyncRegister
  reg_D410
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n705),
    .dout0(n706)
  );


  SyncRegister
  reg_D411
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n688),
    .dout0(n689)
  );


  SyncRegister
  reg_D412
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n706),
    .dout0(n707)
  );


  SyncRegister
  reg_D413
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n689),
    .dout0(n694)
  );


  SyncRegister
  reg_D414
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n707),
    .dout0(n708)
  );


  SyncRegister
  reg_D415
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n708),
    .dout0(n757)
  );


  SyncRegister
  reg_D416
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n698),
    .dout0(n701)
  );


  SyncRegister
  reg_D417
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n712),
    .dout0(n716)
  );


  SyncRegister
  reg_D418
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n720),
    .din0(n756)
  );


  SyncRegister
  reg_D419
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n728),
    .din0(n757)
  );


  SyncRegister
  reg_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n52),
    .dout0(n55)
  );


  SyncRegister
  reg_D420
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n734),
    .din0(n756)
  );


  SyncRegister
  reg_D421
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n728),
    .dout0(n729)
  );


  SyncRegister
  reg_D422
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n720),
    .dout0(n721)
  );


  SyncRegister
  reg_D423
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n721),
    .dout0(n722)
  );


  SyncRegister
  reg_D424
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n729),
    .dout0(n730)
  );


  SyncRegister
  reg_D425
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n722),
    .dout0(n723)
  );


  SyncRegister
  reg_D426
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n730),
    .dout0(n731)
  );


  SyncRegister
  reg_D427
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n723),
    .dout0(n724)
  );


  SyncRegister
  reg_D428
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n724),
    .dout0(n725)
  );


  SyncRegister
  reg_D429
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n742),
    .dout0(n743)
  );


  SyncRegister
  reg_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n66),
    .dout0(n70)
  );


  SyncRegister
  reg_D430
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n742),
    .dout0(n749)
  );


  SyncRegister
  reg_D431
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n725),
    .dout0(n726)
  );


  SyncRegister
  reg_D432
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n743),
    .dout0(n744)
  );


  SyncRegister
  reg_D433
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n726),
    .dout0(n727)
  );


  SyncRegister
  reg_D434
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n744),
    .dout0(n745)
  );


  SyncRegister
  reg_D435
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n727),
    .dout0(n732)
  );


  SyncRegister
  reg_D436
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n745),
    .dout0(n746)
  );


  SyncRegister
  reg_D437
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n746),
    .dout0(n795)
  );


  SyncRegister
  reg_D438
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n736),
    .dout0(n739)
  );


  SyncRegister
  reg_D439
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n750),
    .dout0(n754)
  );


  SyncRegister
  reg_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n110),
    .dout0(n74)
  );


  SyncRegister
  reg_D440
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n758),
    .din0(n794)
  );


  SyncRegister
  reg_D441
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n766),
    .din0(n795)
  );


  SyncRegister
  reg_D442
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n772),
    .din0(n794)
  );


  SyncRegister
  reg_D443
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n766),
    .dout0(n767)
  );


  SyncRegister
  reg_D444
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n758),
    .dout0(n759)
  );


  SyncRegister
  reg_D445
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n759),
    .dout0(n760)
  );


  SyncRegister
  reg_D446
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n767),
    .dout0(n768)
  );


  SyncRegister
  reg_D447
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n760),
    .dout0(n761)
  );


  SyncRegister
  reg_D448
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n768),
    .dout0(n769)
  );


  SyncRegister
  reg_D449
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n761),
    .dout0(n762)
  );


  SyncRegister
  reg_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n111),
    .dout0(n82)
  );


  SyncRegister
  reg_D450
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n762),
    .dout0(n763)
  );


  SyncRegister
  reg_D451
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n780),
    .dout0(n781)
  );


  SyncRegister
  reg_D452
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n780),
    .dout0(n787)
  );


  SyncRegister
  reg_D453
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n763),
    .dout0(n764)
  );


  SyncRegister
  reg_D454
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n781),
    .dout0(n782)
  );


  SyncRegister
  reg_D455
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n764),
    .dout0(n765)
  );


  SyncRegister
  reg_D456
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n782),
    .dout0(n783)
  );


  SyncRegister
  reg_D457
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n765),
    .dout0(n770)
  );


  SyncRegister
  reg_D458
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n783),
    .dout0(n784)
  );


  SyncRegister
  reg_D459
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n784),
    .dout0(n833)
  );


  SyncRegister
  reg_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n110),
    .dout0(n88)
  );


  SyncRegister
  reg_D460
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n774),
    .dout0(n777)
  );


  SyncRegister
  reg_D461
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n788),
    .dout0(n792)
  );


  SyncRegister
  reg_D462
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n796),
    .din0(n832)
  );


  SyncRegister
  reg_D463
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n804),
    .din0(n833)
  );


  SyncRegister
  reg_D464
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n810),
    .din0(n832)
  );


  SyncRegister
  reg_D465
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n804),
    .dout0(n805)
  );


  SyncRegister
  reg_D466
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n796),
    .dout0(n797)
  );


  SyncRegister
  reg_D467
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n797),
    .dout0(n798)
  );


  SyncRegister
  reg_D468
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n805),
    .dout0(n806)
  );


  SyncRegister
  reg_D469
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n798),
    .dout0(n799)
  );


  SyncRegister
  reg_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n82),
    .dout0(n83)
  );


  SyncRegister
  reg_D470
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n806),
    .dout0(n807)
  );


  SyncRegister
  reg_D471
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n799),
    .dout0(n800)
  );


  SyncRegister
  reg_D472
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n800),
    .dout0(n801)
  );


  SyncRegister
  reg_D473
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n818),
    .dout0(n819)
  );


  SyncRegister
  reg_D474
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n818),
    .dout0(n825)
  );


  SyncRegister
  reg_D475
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n801),
    .dout0(n802)
  );


  SyncRegister
  reg_D476
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n819),
    .dout0(n820)
  );


  SyncRegister
  reg_D477
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n802),
    .dout0(n803)
  );


  SyncRegister
  reg_D478
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n820),
    .dout0(n821)
  );


  SyncRegister
  reg_D479
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n803),
    .dout0(n808)
  );


  SyncRegister
  reg_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n74),
    .dout0(n75)
  );


  SyncRegister
  reg_D480
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n821),
    .dout0(n822)
  );


  SyncRegister
  reg_D481
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n822),
    .dout0(n871)
  );


  SyncRegister
  reg_D482
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n812),
    .dout0(n815)
  );


  SyncRegister
  reg_D483
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n826),
    .dout0(n830)
  );


  SyncRegister
  reg_D484
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n834),
    .din0(n870)
  );


  SyncRegister
  reg_D485
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n842),
    .din0(n871)
  );


  SyncRegister
  reg_D486
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n848),
    .din0(n870)
  );


  SyncRegister
  reg_D487
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n842),
    .dout0(n843)
  );


  SyncRegister
  reg_D488
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n834),
    .dout0(n835)
  );


  SyncRegister
  reg_D489
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n835),
    .dout0(n836)
  );


  SyncRegister
  reg_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n75),
    .dout0(n76)
  );


  SyncRegister
  reg_D490
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n843),
    .dout0(n844)
  );


  SyncRegister
  reg_D491
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n836),
    .dout0(n837)
  );


  SyncRegister
  reg_D492
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n844),
    .dout0(n845)
  );


  SyncRegister
  reg_D493
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n837),
    .dout0(n838)
  );


  SyncRegister
  reg_D494
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n838),
    .dout0(n839)
  );


  SyncRegister
  reg_D495
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n856),
    .dout0(n857)
  );


  SyncRegister
  reg_D496
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n856),
    .dout0(n863)
  );


  SyncRegister
  reg_D497
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n839),
    .dout0(n840)
  );


  SyncRegister
  reg_D498
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n857),
    .dout0(n858)
  );


  SyncRegister
  reg_D499
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n840),
    .dout0(n841)
  );


  SyncRegister
  reg_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1),
    .dout0(n2)
  );


  SyncRegister
  reg_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n83),
    .dout0(n84)
  );


  SyncRegister
  reg_D500
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n858),
    .dout0(n859)
  );


  SyncRegister
  reg_D501
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n841),
    .dout0(n846)
  );


  SyncRegister
  reg_D502
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n859),
    .dout0(n860)
  );


  SyncRegister
  reg_D503
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n860),
    .dout0(n909)
  );


  SyncRegister
  reg_D504
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n850),
    .dout0(n853)
  );


  SyncRegister
  reg_D505
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n864),
    .dout0(n868)
  );


  SyncRegister
  reg_D506
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n872),
    .din0(n908)
  );


  SyncRegister
  reg_D507
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n880),
    .din0(n909)
  );


  SyncRegister
  reg_D508
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n886),
    .din0(n908)
  );


  SyncRegister
  reg_D509
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n880),
    .dout0(n881)
  );


  SyncRegister
  reg_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n76),
    .dout0(n77)
  );


  SyncRegister
  reg_D510
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n872),
    .dout0(n873)
  );


  SyncRegister
  reg_D511
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n873),
    .dout0(n874)
  );


  SyncRegister
  reg_D512
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n881),
    .dout0(n882)
  );


  SyncRegister
  reg_D513
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n874),
    .dout0(n875)
  );


  SyncRegister
  reg_D514
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n882),
    .dout0(n883)
  );


  SyncRegister
  reg_D515
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n875),
    .dout0(n876)
  );


  SyncRegister
  reg_D516
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n876),
    .dout0(n877)
  );


  SyncRegister
  reg_D517
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n894),
    .dout0(n895)
  );


  SyncRegister
  reg_D518
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n894),
    .dout0(n901)
  );


  SyncRegister
  reg_D519
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n877),
    .dout0(n878)
  );


  SyncRegister
  reg_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n84),
    .dout0(n85)
  );


  SyncRegister
  reg_D520
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n895),
    .dout0(n896)
  );


  SyncRegister
  reg_D521
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n878),
    .dout0(n879)
  );


  SyncRegister
  reg_D522
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n896),
    .dout0(n897)
  );


  SyncRegister
  reg_D523
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n879),
    .dout0(n884)
  );


  SyncRegister
  reg_D524
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n897),
    .dout0(n898)
  );


  SyncRegister
  reg_D525
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n898),
    .dout0(n947)
  );


  SyncRegister
  reg_D526
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n888),
    .dout0(n891)
  );


  SyncRegister
  reg_D527
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n902),
    .dout0(n906)
  );


  SyncRegister
  reg_D528
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n910),
    .din0(n946)
  );


  SyncRegister
  reg_D529
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n918),
    .din0(n947)
  );


  SyncRegister
  reg_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n77),
    .dout0(n78)
  );


  SyncRegister
  reg_D530
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n924),
    .din0(n946)
  );


  SyncRegister
  reg_D531
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n918),
    .dout0(n919)
  );


  SyncRegister
  reg_D532
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n910),
    .dout0(n911)
  );


  SyncRegister
  reg_D533
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n911),
    .dout0(n912)
  );


  SyncRegister
  reg_D534
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n919),
    .dout0(n920)
  );


  SyncRegister
  reg_D535
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n912),
    .dout0(n913)
  );


  SyncRegister
  reg_D536
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n920),
    .dout0(n921)
  );


  SyncRegister
  reg_D537
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n913),
    .dout0(n914)
  );


  SyncRegister
  reg_D538
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n914),
    .dout0(n915)
  );


  SyncRegister
  reg_D539
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n932),
    .dout0(n933)
  );


  SyncRegister
  reg_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n78),
    .dout0(n79)
  );


  SyncRegister
  reg_D540
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n932),
    .dout0(n939)
  );


  SyncRegister
  reg_D541
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n915),
    .dout0(n916)
  );


  SyncRegister
  reg_D542
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n933),
    .dout0(n934)
  );


  SyncRegister
  reg_D543
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n916),
    .dout0(n917)
  );


  SyncRegister
  reg_D544
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n934),
    .dout0(n935)
  );


  SyncRegister
  reg_D545
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n917),
    .dout0(n922)
  );


  SyncRegister
  reg_D546
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n935),
    .dout0(n936)
  );


  SyncRegister
  reg_D547
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n936),
    .dout0(n985)
  );


  SyncRegister
  reg_D548
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n926),
    .dout0(n929)
  );


  SyncRegister
  reg_D549
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n940),
    .dout0(n944)
  );


  SyncRegister
  reg_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n96),
    .dout0(n97)
  );


  SyncRegister
  reg_D550
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n948),
    .din0(n984)
  );


  SyncRegister
  reg_D551
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n956),
    .din0(n985)
  );


  SyncRegister
  reg_D552
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n962),
    .din0(n984)
  );


  SyncRegister
  reg_D553
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n956),
    .dout0(n957)
  );


  SyncRegister
  reg_D554
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n948),
    .dout0(n949)
  );


  SyncRegister
  reg_D555
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n949),
    .dout0(n950)
  );


  SyncRegister
  reg_D556
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n957),
    .dout0(n958)
  );


  SyncRegister
  reg_D557
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n950),
    .dout0(n951)
  );


  SyncRegister
  reg_D558
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n958),
    .dout0(n959)
  );


  SyncRegister
  reg_D559
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n951),
    .dout0(n952)
  );


  SyncRegister
  reg_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n103),
    .din0(n96)
  );


  SyncRegister
  reg_D560
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n952),
    .dout0(n953)
  );


  SyncRegister
  reg_D561
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n970),
    .dout0(n971)
  );


  SyncRegister
  reg_D562
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n970),
    .dout0(n977)
  );


  SyncRegister
  reg_D563
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n953),
    .dout0(n954)
  );


  SyncRegister
  reg_D564
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n971),
    .dout0(n972)
  );


  SyncRegister
  reg_D565
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n954),
    .dout0(n955)
  );


  SyncRegister
  reg_D566
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n972),
    .dout0(n973)
  );


  SyncRegister
  reg_D567
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n955),
    .dout0(n960)
  );


  SyncRegister
  reg_D568
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n973),
    .dout0(n974)
  );


  SyncRegister
  reg_D569
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1023),
    .din0(n974)
  );


  SyncRegister
  reg_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n79),
    .dout0(n80)
  );


  SyncRegister
  reg_D570
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n964),
    .dout0(n967)
  );


  SyncRegister
  reg_D571
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n978),
    .dout0(n982)
  );


  SyncRegister
  reg_D572
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1022),
    .dout0(n986)
  );


  SyncRegister
  reg_D573
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1023),
    .dout0(n994)
  );


  SyncRegister
  reg_D574
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1000),
    .din0(n1022)
  );


  SyncRegister
  reg_D575
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n994),
    .dout0(n995)
  );


  SyncRegister
  reg_D576
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n986),
    .dout0(n987)
  );


  SyncRegister
  reg_D577
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n987),
    .dout0(n988)
  );


  SyncRegister
  reg_D578
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n995),
    .dout0(n996)
  );


  SyncRegister
  reg_D579
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n988),
    .dout0(n989)
  );


  SyncRegister
  reg_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n97),
    .dout0(n98)
  );


  SyncRegister
  reg_D580
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n996),
    .dout0(n997)
  );


  SyncRegister
  reg_D581
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n989),
    .dout0(n990)
  );


  SyncRegister
  reg_D582
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n990),
    .dout0(n991)
  );


  SyncRegister
  reg_D583
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1008),
    .dout0(n1009)
  );


  SyncRegister
  reg_D584
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1008),
    .dout0(n1015)
  );


  SyncRegister
  reg_D585
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n991),
    .dout0(n992)
  );


  SyncRegister
  reg_D586
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1009),
    .dout0(n1010)
  );


  SyncRegister
  reg_D587
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n992),
    .dout0(n993)
  );


  SyncRegister
  reg_D588
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1010),
    .dout0(n1011)
  );


  SyncRegister
  reg_D589
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n993),
    .dout0(n998)
  );


  SyncRegister
  reg_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n80),
    .dout0(n81)
  );


  SyncRegister
  reg_D590
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1011),
    .dout0(n1012)
  );


  SyncRegister
  reg_D591
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1012),
    .dout0(n1061)
  );


  SyncRegister
  reg_D592
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1002),
    .dout0(n1005)
  );


  SyncRegister
  reg_D593
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1016),
    .dout0(n1020)
  );


  SyncRegister
  reg_D594
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1024),
    .din0(n1060)
  );


  SyncRegister
  reg_D595
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1032),
    .din0(n1061)
  );


  SyncRegister
  reg_D596
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1038),
    .din0(n1060)
  );


  SyncRegister
  reg_D597
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1032),
    .dout0(n1033)
  );


  SyncRegister
  reg_D598
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1024),
    .dout0(n1025)
  );


  SyncRegister
  reg_D599
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1025),
    .dout0(n1026)
  );


  SyncRegister
  reg_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n10),
    .din0(n9)
  );


  SyncRegister
  reg_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n98),
    .dout0(n99)
  );


  SyncRegister
  reg_D600
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1033),
    .dout0(n1034)
  );


  SyncRegister
  reg_D601
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1026),
    .dout0(n1027)
  );


  SyncRegister
  reg_D602
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1034),
    .dout0(n1035)
  );


  SyncRegister
  reg_D603
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1027),
    .dout0(n1028)
  );


  SyncRegister
  reg_D604
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1028),
    .dout0(n1029)
  );


  SyncRegister
  reg_D605
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1046),
    .dout0(n1047)
  );


  SyncRegister
  reg_D606
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1046),
    .dout0(n1053)
  );


  SyncRegister
  reg_D607
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1029),
    .dout0(n1030)
  );


  SyncRegister
  reg_D608
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1047),
    .dout0(n1048)
  );


  SyncRegister
  reg_D609
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1030),
    .dout0(n1031)
  );


  SyncRegister
  reg_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n81),
    .dout0(n86)
  );


  SyncRegister
  reg_D610
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1048),
    .dout0(n1049)
  );


  SyncRegister
  reg_D611
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1031),
    .dout0(n1036)
  );


  SyncRegister
  reg_D612
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1049),
    .dout0(n1050)
  );


  SyncRegister
  reg_D613
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1050),
    .dout0(n1099)
  );


  SyncRegister
  reg_D614
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1040),
    .dout0(n1043)
  );


  SyncRegister
  reg_D615
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1054),
    .dout0(n1058)
  );


  SyncRegister
  reg_D616
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1062),
    .din0(n1098)
  );


  SyncRegister
  reg_D617
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1070),
    .din0(n1099)
  );


  SyncRegister
  reg_D618
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1076),
    .din0(n1098)
  );


  SyncRegister
  reg_D619
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1070),
    .dout0(n1071)
  );


  SyncRegister
  reg_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n100),
    .din0(n99)
  );


  SyncRegister
  reg_D620
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1062),
    .dout0(n1063)
  );


  SyncRegister
  reg_D621
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1063),
    .dout0(n1064)
  );


  SyncRegister
  reg_D622
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1071),
    .dout0(n1072)
  );


  SyncRegister
  reg_D623
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1064),
    .dout0(n1065)
  );


  SyncRegister
  reg_D624
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1072),
    .dout0(n1073)
  );


  SyncRegister
  reg_D625
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1065),
    .dout0(n1066)
  );


  SyncRegister
  reg_D626
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1066),
    .dout0(n1067)
  );


  SyncRegister
  reg_D627
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1084),
    .dout0(n1085)
  );


  SyncRegister
  reg_D628
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1084),
    .dout0(n1091)
  );


  SyncRegister
  reg_D629
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1067),
    .dout0(n1068)
  );


  SyncRegister
  reg_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n100),
    .dout0(n149)
  );


  SyncRegister
  reg_D630
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1085),
    .dout0(n1086)
  );


  SyncRegister
  reg_D631
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1068),
    .dout0(n1069)
  );


  SyncRegister
  reg_D632
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1086),
    .dout0(n1087)
  );


  SyncRegister
  reg_D633
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1069),
    .dout0(n1074)
  );


  SyncRegister
  reg_D634
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1087),
    .dout0(n1088)
  );


  SyncRegister
  reg_D635
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1088),
    .dout0(n1137)
  );


  SyncRegister
  reg_D636
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1078),
    .dout0(n1081)
  );


  SyncRegister
  reg_D637
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1092),
    .dout0(n1096)
  );


  SyncRegister
  reg_D638
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1100),
    .din0(n1136)
  );


  SyncRegister
  reg_D639
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1108),
    .din0(n1137)
  );


  SyncRegister
  reg_D64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n90),
    .dout0(n93)
  );


  SyncRegister
  reg_D640
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1114),
    .din0(n1136)
  );


  SyncRegister
  reg_D641
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1108),
    .dout0(n1109)
  );


  SyncRegister
  reg_D642
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1100),
    .dout0(n1101)
  );


  SyncRegister
  reg_D643
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1101),
    .dout0(n1102)
  );


  SyncRegister
  reg_D644
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1109),
    .dout0(n1110)
  );


  SyncRegister
  reg_D645
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1102),
    .dout0(n1103)
  );


  SyncRegister
  reg_D646
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1110),
    .dout0(n1111)
  );


  SyncRegister
  reg_D647
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1103),
    .dout0(n1104)
  );


  SyncRegister
  reg_D648
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1104),
    .dout0(n1105)
  );


  SyncRegister
  reg_D649
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1122),
    .dout0(n1123)
  );


  SyncRegister
  reg_D65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n104),
    .dout0(n108)
  );


  SyncRegister
  reg_D650
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1122),
    .dout0(n1129)
  );


  SyncRegister
  reg_D651
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1105),
    .dout0(n1106)
  );


  SyncRegister
  reg_D652
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1123),
    .dout0(n1124)
  );


  SyncRegister
  reg_D653
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1106),
    .dout0(n1107)
  );


  SyncRegister
  reg_D654
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1124),
    .dout0(n1125)
  );


  SyncRegister
  reg_D655
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1107),
    .dout0(n1112)
  );


  SyncRegister
  reg_D656
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1125),
    .dout0(n1126)
  );


  SyncRegister
  reg_D657
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1126),
    .dout0(n1175)
  );


  SyncRegister
  reg_D658
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1116),
    .dout0(n1119)
  );


  SyncRegister
  reg_D659
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1130),
    .dout0(n1134)
  );


  SyncRegister
  reg_D66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n112),
    .din0(n148)
  );


  SyncRegister
  reg_D660
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1138),
    .din0(n1174)
  );


  SyncRegister
  reg_D661
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1146),
    .din0(n1175)
  );


  SyncRegister
  reg_D662
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1152),
    .din0(n1174)
  );


  SyncRegister
  reg_D663
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1146),
    .dout0(n1147)
  );


  SyncRegister
  reg_D664
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1138),
    .dout0(n1139)
  );


  SyncRegister
  reg_D665
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1139),
    .dout0(n1140)
  );


  SyncRegister
  reg_D666
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1147),
    .dout0(n1148)
  );


  SyncRegister
  reg_D667
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1140),
    .dout0(n1141)
  );


  SyncRegister
  reg_D668
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1148),
    .dout0(n1149)
  );


  SyncRegister
  reg_D669
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1141),
    .dout0(n1142)
  );


  SyncRegister
  reg_D67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n120),
    .din0(n149)
  );


  SyncRegister
  reg_D670
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1142),
    .dout0(n1143)
  );


  SyncRegister
  reg_D671
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1160),
    .dout0(n1161)
  );


  SyncRegister
  reg_D672
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1160),
    .dout0(n1167)
  );


  SyncRegister
  reg_D673
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1143),
    .dout0(n1144)
  );


  SyncRegister
  reg_D674
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1161),
    .dout0(n1162)
  );


  SyncRegister
  reg_D675
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1144),
    .dout0(n1145)
  );


  SyncRegister
  reg_D676
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1162),
    .dout0(n1163)
  );


  SyncRegister
  reg_D677
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1145),
    .dout0(n1150)
  );


  SyncRegister
  reg_D678
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1163),
    .dout0(n1164)
  );


  SyncRegister
  reg_D679
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1164),
    .dout0(n1213)
  );


  SyncRegister
  reg_D68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n126),
    .din0(n148)
  );


  SyncRegister
  reg_D680
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1154),
    .dout0(n1157)
  );


  SyncRegister
  reg_D681
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1168),
    .dout0(n1172)
  );


  SyncRegister
  reg_D682
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1176),
    .din0(n1212)
  );


  SyncRegister
  reg_D683
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1184),
    .din0(n1213)
  );


  SyncRegister
  reg_D684
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1190),
    .din0(n1212)
  );


  SyncRegister
  reg_D685
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1184),
    .dout0(n1185)
  );


  SyncRegister
  reg_D686
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1176),
    .dout0(n1177)
  );


  SyncRegister
  reg_D687
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1177),
    .dout0(n1178)
  );


  SyncRegister
  reg_D688
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1185),
    .dout0(n1186)
  );


  SyncRegister
  reg_D689
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1178),
    .dout0(n1179)
  );


  SyncRegister
  reg_D69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n120),
    .dout0(n121)
  );


  SyncRegister
  reg_D690
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1186),
    .dout0(n1187)
  );


  SyncRegister
  reg_D691
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1179),
    .dout0(n1180)
  );


  SyncRegister
  reg_D692
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1180),
    .dout0(n1181)
  );


  SyncRegister
  reg_D693
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1198),
    .dout0(n1199)
  );


  SyncRegister
  reg_D694
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1198),
    .dout0(n1205)
  );


  SyncRegister
  reg_D695
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1181),
    .dout0(n1182)
  );


  SyncRegister
  reg_D696
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1199),
    .dout0(n1200)
  );


  SyncRegister
  reg_D697
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1182),
    .dout0(n1183)
  );


  SyncRegister
  reg_D698
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1200),
    .dout0(n1201)
  );


  SyncRegister
  reg_D699
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1183),
    .dout0(n1188)
  );


  SyncRegister
  reg_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2),
    .dout0(n3)
  );


  SyncRegister
  reg_D70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n112),
    .dout0(n113)
  );


  SyncRegister
  reg_D700
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1201),
    .dout0(n1202)
  );


  SyncRegister
  reg_D701
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1202),
    .dout0(n1215)
  );


  SyncRegister
  reg_D702
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1192),
    .dout0(n1195)
  );


  SyncRegister
  reg_D703
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1206),
    .dout0(n1210)
  );


  SyncRegister
  reg_D71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n113),
    .dout0(n114)
  );


  SyncRegister
  reg_D72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n121),
    .dout0(n122)
  );


  SyncRegister
  reg_D73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n114),
    .dout0(n115)
  );


  SyncRegister
  reg_D74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n122),
    .dout0(n123)
  );


  SyncRegister
  reg_D75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n115),
    .dout0(n116)
  );


  SyncRegister
  reg_D76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n116),
    .dout0(n117)
  );


  SyncRegister
  reg_D77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n134),
    .dout0(n135)
  );


  SyncRegister
  reg_D78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n134),
    .dout0(n141)
  );


  SyncRegister
  reg_D79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n117),
    .dout0(n118)
  );


  SyncRegister
  reg_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n10),
    .dout0(n11)
  );


  SyncRegister
  reg_D80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n135),
    .dout0(n136)
  );


  SyncRegister
  reg_D81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n118),
    .dout0(n119)
  );


  SyncRegister
  reg_D82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n136),
    .dout0(n137)
  );


  SyncRegister
  reg_D83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n119),
    .dout0(n124)
  );


  SyncRegister
  reg_D84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n137),
    .dout0(n138)
  );


  SyncRegister
  reg_D85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n138),
    .dout0(n187)
  );


  SyncRegister
  reg_D86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n128),
    .dout0(n131)
  );


  SyncRegister
  reg_D87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n142),
    .dout0(n146)
  );


  SyncRegister
  reg_D88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n150),
    .din0(n186)
  );


  SyncRegister
  reg_D89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n158),
    .din0(n187)
  );


  SyncRegister
  reg_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n3),
    .dout0(n4)
  );


  SyncRegister
  reg_D90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n164),
    .din0(n186)
  );


  SyncRegister
  reg_D91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n158),
    .dout0(n159)
  );


  SyncRegister
  reg_D92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n150),
    .dout0(n151)
  );


  SyncRegister
  reg_D93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n151),
    .dout0(n152)
  );


  SyncRegister
  reg_D94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n159),
    .dout0(n160)
  );


  SyncRegister
  reg_D95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n152),
    .dout0(n153)
  );


  SyncRegister
  reg_D96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n160),
    .dout0(n161)
  );


  SyncRegister
  reg_D97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n153),
    .dout0(n154)
  );


  SyncRegister
  reg_D98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n154),
    .dout0(n155)
  );


  SyncRegister
  reg_D99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n172),
    .dout0(n173)
  );


  SyncRegister
  reg_fir0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1216),
    .dout0(n1218)
  );


  SyncRegister
  reg_fir1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1217),
    .dout0(n1219)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1243),
    .din0(n2446)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1252),
    .dout0(n1257)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1431),
    .din0(n1454)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1440),
    .dout0(n1445)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1469),
    .din0(n1492)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1478),
    .dout0(n1483)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1507),
    .din0(n1530)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1516),
    .dout0(n1521)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1545),
    .din0(n1568)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1554),
    .dout0(n1559)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1583),
    .din0(n1606)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1592),
    .dout0(n1597)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1279),
    .din0(n1302)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1621),
    .din0(n1644)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1630),
    .dout0(n1635)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1659),
    .din0(n1682)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1668),
    .dout0(n1673)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1697),
    .din0(n1720)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1706),
    .dout0(n1711)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1735),
    .din0(n1758)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1744),
    .dout0(n1749)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1773),
    .din0(n1796)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1782),
    .dout0(n1787)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1288),
    .dout0(n1293)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1811),
    .din0(n1834)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1820),
    .dout0(n1825)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1849),
    .din0(n1872)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1858),
    .dout0(n1863)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1887),
    .din0(n1910)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1896),
    .dout0(n1901)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1925),
    .din0(n1948)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1934),
    .dout0(n1939)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1963),
    .din0(n1986)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1972),
    .dout0(n1977)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1317),
    .din0(n1340)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2001),
    .din0(n2024)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2010),
    .dout0(n2015)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2039),
    .din0(n2062)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2048),
    .dout0(n2053)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2077),
    .din0(n2100)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2086),
    .dout0(n2091)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2115),
    .din0(n2138)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2124),
    .dout0(n2129)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2153),
    .din0(n2176)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2162),
    .dout0(n2167)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1326),
    .dout0(n1331)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2191),
    .din0(n2214)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2200),
    .dout0(n2205)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2229),
    .din0(n2252)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2238),
    .dout0(n2243)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2267),
    .din0(n2290)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2276),
    .dout0(n2281)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2305),
    .din0(n2328)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2314),
    .dout0(n2319)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2343),
    .din0(n2366)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2352),
    .dout0(n2357)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1355),
    .din0(n1378)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2381),
    .din0(n2404)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2390),
    .dout0(n2395)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2419),
    .din0(n2442)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2428),
    .dout0(n2433)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1364),
    .dout0(n1369)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1393),
    .din0(n1416)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1402),
    .dout0(n1407)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n13),
    .din0(n2444)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n22),
    .dout0(n27)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n201),
    .din0(n224)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n210),
    .dout0(n215)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n239),
    .din0(n262)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n248),
    .dout0(n253)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n277),
    .din0(n300)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n286),
    .dout0(n291)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n315),
    .din0(n338)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n324),
    .dout0(n329)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n353),
    .din0(n376)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n362),
    .dout0(n367)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n49),
    .din0(n72)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n391),
    .din0(n414)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n400),
    .dout0(n405)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n429),
    .din0(n452)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n438),
    .dout0(n443)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n467),
    .din0(n490)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n476),
    .dout0(n481)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n505),
    .din0(n528)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n514),
    .dout0(n519)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n543),
    .din0(n566)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n552),
    .dout0(n557)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n58),
    .dout0(n63)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n581),
    .din0(n604)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n590),
    .dout0(n595)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n619),
    .din0(n642)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n628),
    .dout0(n633)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n657),
    .din0(n680)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n666),
    .dout0(n671)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n695),
    .din0(n718)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n704),
    .dout0(n709)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n733),
    .din0(n756)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n742),
    .dout0(n747)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n110),
    .dout0(n87)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n771),
    .din0(n794)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n780),
    .dout0(n785)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n809),
    .din0(n832)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n818),
    .dout0(n823)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n847),
    .din0(n870)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n856),
    .dout0(n861)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n885),
    .din0(n908)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n894),
    .dout0(n899)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n923),
    .din0(n946)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n932),
    .dout0(n937)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n101),
    .din0(n96)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n961),
    .din0(n984)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n970),
    .dout0(n975)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1022),
    .dout0(n999)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1008),
    .dout0(n1013)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1037),
    .din0(n1060)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1046),
    .dout0(n1051)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1075),
    .din0(n1098)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1084),
    .dout0(n1089)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1113),
    .din0(n1136)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1122),
    .dout0(n1127)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n125),
    .din0(n148)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1151),
    .din0(n1174)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1160),
    .dout0(n1165)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1189),
    .din0(n1212)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1198),
    .dout0(n1203)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n134),
    .dout0(n139)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n163),
    .din0(n186)
  );


  SyncShlI
  #(
    .ID(1),
    .IMMEDIATE(4)
  )
  shli_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n172),
    .dout0(n177)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1245),
    .din0(n2446)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1252),
    .dout0(n1258)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1433),
    .din0(n1454)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1440),
    .dout0(n1446)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1471),
    .din0(n1492)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1478),
    .dout0(n1484)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1509),
    .din0(n1530)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1516),
    .dout0(n1522)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1547),
    .din0(n1568)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1554),
    .dout0(n1560)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1585),
    .din0(n1606)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1592),
    .dout0(n1598)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1281),
    .din0(n1302)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1623),
    .din0(n1644)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1630),
    .dout0(n1636)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1661),
    .din0(n1682)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1668),
    .dout0(n1674)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1699),
    .din0(n1720)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1706),
    .dout0(n1712)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1737),
    .din0(n1758)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1744),
    .dout0(n1750)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1775),
    .din0(n1796)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1782),
    .dout0(n1788)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1288),
    .dout0(n1294)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1813),
    .din0(n1834)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1820),
    .dout0(n1826)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1851),
    .din0(n1872)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1858),
    .dout0(n1864)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1889),
    .din0(n1910)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1896),
    .dout0(n1902)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1927),
    .din0(n1948)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1934),
    .dout0(n1940)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1965),
    .din0(n1986)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1972),
    .dout0(n1978)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1319),
    .din0(n1340)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2003),
    .din0(n2024)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2010),
    .dout0(n2016)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2041),
    .din0(n2062)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2048),
    .dout0(n2054)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2079),
    .din0(n2100)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2086),
    .dout0(n2092)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2117),
    .din0(n2138)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2124),
    .dout0(n2130)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2155),
    .din0(n2176)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2162),
    .dout0(n2168)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1326),
    .dout0(n1332)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2193),
    .din0(n2214)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2200),
    .dout0(n2206)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2231),
    .din0(n2252)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2238),
    .dout0(n2244)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2269),
    .din0(n2290)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2276),
    .dout0(n2282)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2307),
    .din0(n2328)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2314),
    .dout0(n2320)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2345),
    .din0(n2366)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2352),
    .dout0(n2358)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1357),
    .din0(n1378)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2383),
    .din0(n2404)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2390),
    .dout0(n2396)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n2421),
    .din0(n2442)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2428),
    .dout0(n2434)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1364),
    .dout0(n1370)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1395),
    .din0(n1416)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1402),
    .dout0(n1408)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n15),
    .din0(n2444)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n22),
    .dout0(n28)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n203),
    .din0(n224)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n210),
    .dout0(n216)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n241),
    .din0(n262)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n248),
    .dout0(n254)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n279),
    .din0(n300)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n286),
    .dout0(n292)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n317),
    .din0(n338)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n324),
    .dout0(n330)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n355),
    .din0(n376)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n362),
    .dout0(n368)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n51),
    .din0(n72)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n393),
    .din0(n414)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n400),
    .dout0(n406)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n431),
    .din0(n452)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n438),
    .dout0(n444)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n469),
    .din0(n490)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n476),
    .dout0(n482)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n507),
    .din0(n528)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n514),
    .dout0(n520)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n545),
    .din0(n566)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n552),
    .dout0(n558)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n58),
    .dout0(n64)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n583),
    .din0(n604)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n590),
    .dout0(n596)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n621),
    .din0(n642)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n628),
    .dout0(n634)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n659),
    .din0(n680)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n666),
    .dout0(n672)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n697),
    .din0(n718)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n704),
    .dout0(n710)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n735),
    .din0(n756)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n742),
    .dout0(n748)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n110),
    .dout0(n89)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n773),
    .din0(n794)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n780),
    .dout0(n786)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n811),
    .din0(n832)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n818),
    .dout0(n824)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n849),
    .din0(n870)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n856),
    .dout0(n862)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n887),
    .din0(n908)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n894),
    .dout0(n900)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n925),
    .din0(n946)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n932),
    .dout0(n938)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n102),
    .din0(n96)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n963),
    .din0(n984)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n970),
    .dout0(n976)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1001),
    .din0(n1022)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1008),
    .dout0(n1014)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1039),
    .din0(n1060)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1046),
    .dout0(n1052)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1077),
    .din0(n1098)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1084),
    .dout0(n1090)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1115),
    .din0(n1136)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1122),
    .dout0(n1128)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n127),
    .din0(n148)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1153),
    .din0(n1174)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1160),
    .dout0(n1166)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1191),
    .din0(n1212)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1198),
    .dout0(n1204)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n134),
    .dout0(n140)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n165),
    .din0(n186)
  );


  SyncShrI
  #(
    .ID(1),
    .IMMEDIATE(5)
  )
  shri_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n172),
    .dout0(n178)
  );


  SyncSub
  sub_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n12),
    .din1(n35),
    .dout0(n72)
  );


  SyncSub
  sub_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n11),
    .din1(n21),
    .dout0(n22)
  );


  SyncSub
  sub_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n200),
    .din1(n223),
    .dout0(n262)
  );


  SyncSub
  sub_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n199),
    .din1(n209),
    .dout0(n210)
  );


  SyncSub
  sub_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n238),
    .din1(n261),
    .dout0(n300)
  );


  SyncSub
  sub_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n237),
    .din1(n247),
    .dout0(n248)
  );


  SyncSub
  sub_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n276),
    .din1(n299),
    .dout0(n338)
  );


  SyncSub
  sub_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n275),
    .din1(n285),
    .dout0(n286)
  );


  SyncSub
  sub_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n314),
    .din1(n337),
    .dout0(n376)
  );


  SyncSub
  sub_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n313),
    .din1(n323),
    .dout0(n324)
  );


  SyncSub
  sub_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n352),
    .din1(n375),
    .dout0(n414)
  );


  SyncSub
  sub_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n351),
    .din1(n361),
    .dout0(n362)
  );


  SyncSub
  sub_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n110),
    .din0(n48),
    .din1(n71)
  );


  SyncSub
  sub_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n390),
    .din1(n413),
    .dout0(n452)
  );


  SyncSub
  sub_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n389),
    .din1(n399),
    .dout0(n400)
  );


  SyncSub
  sub_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n428),
    .din1(n451),
    .dout0(n490)
  );


  SyncSub
  sub_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n427),
    .din1(n437),
    .dout0(n438)
  );


  SyncSub
  sub_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n466),
    .din1(n489),
    .dout0(n528)
  );


  SyncSub
  sub_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n465),
    .din1(n475),
    .dout0(n476)
  );


  SyncSub
  sub_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n504),
    .din1(n527),
    .dout0(n566)
  );


  SyncSub
  sub_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n503),
    .din1(n513),
    .dout0(n514)
  );


  SyncSub
  sub_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n542),
    .din1(n565),
    .dout0(n604)
  );


  SyncSub
  sub_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n541),
    .din1(n551),
    .dout0(n552)
  );


  SyncSub
  sub_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n47),
    .din1(n57),
    .dout0(n58)
  );


  SyncSub
  sub_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n580),
    .din1(n603),
    .dout0(n642)
  );


  SyncSub
  sub_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n579),
    .din1(n589),
    .dout0(n590)
  );


  SyncSub
  sub_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n618),
    .din1(n641),
    .dout0(n680)
  );


  SyncSub
  sub_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n617),
    .din1(n627),
    .dout0(n628)
  );


  SyncSub
  sub_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n656),
    .din1(n679),
    .dout0(n718)
  );


  SyncSub
  sub_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n655),
    .din1(n665),
    .dout0(n666)
  );


  SyncSub
  sub_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n694),
    .din1(n717),
    .dout0(n756)
  );


  SyncSub
  sub_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n693),
    .din1(n703),
    .dout0(n704)
  );


  SyncSub
  sub_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n732),
    .din1(n755),
    .dout0(n794)
  );


  SyncSub
  sub_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n731),
    .din1(n741),
    .dout0(n742)
  );


  SyncSub
  sub_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n109),
    .dout0(n148),
    .din0(n86)
  );


  SyncSub
  sub_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n770),
    .din1(n793),
    .dout0(n832)
  );


  SyncSub
  sub_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n769),
    .din1(n779),
    .dout0(n780)
  );


  SyncSub
  sub_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n808),
    .din1(n831),
    .dout0(n870)
  );


  SyncSub
  sub_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n807),
    .din1(n817),
    .dout0(n818)
  );


  SyncSub
  sub_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n846),
    .din1(n869),
    .dout0(n908)
  );


  SyncSub
  sub_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n845),
    .din1(n855),
    .dout0(n856)
  );


  SyncSub
  sub_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n884),
    .din1(n907),
    .dout0(n946)
  );


  SyncSub
  sub_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n883),
    .din1(n893),
    .dout0(n894)
  );


  SyncSub
  sub_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n922),
    .din1(n945),
    .dout0(n984)
  );


  SyncSub
  sub_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n921),
    .din1(n931),
    .dout0(n932)
  );


  SyncSub
  sub_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n85),
    .din1(n95),
    .dout0(n96)
  );


  SyncSub
  sub_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .dout0(n1022),
    .din0(n960),
    .din1(n983)
  );


  SyncSub
  sub_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n959),
    .din1(n969),
    .dout0(n970)
  );


  SyncSub
  sub_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1021),
    .dout0(n1060),
    .din0(n998)
  );


  SyncSub
  sub_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1007),
    .dout0(n1008),
    .din0(n997)
  );


  SyncSub
  sub_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1036),
    .din1(n1059),
    .dout0(n1098)
  );


  SyncSub
  sub_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1035),
    .din1(n1045),
    .dout0(n1046)
  );


  SyncSub
  sub_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1074),
    .din1(n1097),
    .dout0(n1136)
  );


  SyncSub
  sub_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1073),
    .din1(n1083),
    .dout0(n1084)
  );


  SyncSub
  sub_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1112),
    .din1(n1135),
    .dout0(n1174)
  );


  SyncSub
  sub_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1111),
    .din1(n1121),
    .dout0(n1122)
  );


  SyncSub
  sub_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n124),
    .din1(n147),
    .dout0(n186)
  );


  SyncSub
  sub_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1150),
    .din1(n1173),
    .dout0(n1212)
  );


  SyncSub
  sub_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1149),
    .din1(n1159),
    .dout0(n1160)
  );


  SyncSub
  sub_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1188),
    .din1(n1211),
    .dout0(n1214)
  );


  SyncSub
  sub_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1187),
    .din1(n1197),
    .dout0(n1198)
  );


  SyncSub
  sub_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n123),
    .din1(n133),
    .dout0(n134)
  );


  SyncSub
  sub_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n162),
    .din1(n185),
    .dout0(n224)
  );


  SyncSub
  sub_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n161),
    .din1(n171),
    .dout0(n172)
  );


  SyncXor
  xor_C0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1247),
    .din0(n1248),
    .dout0(n1250)
  );


  SyncXor
  xor_C1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1249),
    .din0(n1250),
    .dout0(n1251)
  );


  SyncXor
  xor_C10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1335),
    .din1(n1336),
    .dout0(n1337)
  );


  SyncXor
  xor_C100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2195),
    .din0(n2196),
    .dout0(n2198)
  );


  SyncXor
  xor_C101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2197),
    .din0(n2198),
    .dout0(n2199)
  );


  SyncXor
  xor_C102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2209),
    .din1(n2210),
    .dout0(n2211)
  );


  SyncXor
  xor_C103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2211),
    .din1(n2212),
    .dout0(n2213)
  );


  SyncXor
  xor_C104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2233),
    .din0(n2234),
    .dout0(n2236)
  );


  SyncXor
  xor_C105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2235),
    .din0(n2236),
    .dout0(n2237)
  );


  SyncXor
  xor_C106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2247),
    .din1(n2248),
    .dout0(n2249)
  );


  SyncXor
  xor_C107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2249),
    .din1(n2250),
    .dout0(n2251)
  );


  SyncXor
  xor_C108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2271),
    .din0(n2272),
    .dout0(n2274)
  );


  SyncXor
  xor_C109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2273),
    .din0(n2274),
    .dout0(n2275)
  );


  SyncXor
  xor_C11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1337),
    .din1(n1338),
    .dout0(n1339)
  );


  SyncXor
  xor_C110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2285),
    .din1(n2286),
    .dout0(n2287)
  );


  SyncXor
  xor_C111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2287),
    .din1(n2288),
    .dout0(n2289)
  );


  SyncXor
  xor_C112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2309),
    .din0(n2310),
    .dout0(n2312)
  );


  SyncXor
  xor_C113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2311),
    .din0(n2312),
    .dout0(n2313)
  );


  SyncXor
  xor_C114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2323),
    .din1(n2324),
    .dout0(n2325)
  );


  SyncXor
  xor_C115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2325),
    .din1(n2326),
    .dout0(n2327)
  );


  SyncXor
  xor_C116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2347),
    .din0(n2348),
    .dout0(n2350)
  );


  SyncXor
  xor_C117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2349),
    .din0(n2350),
    .dout0(n2351)
  );


  SyncXor
  xor_C118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2361),
    .din1(n2362),
    .dout0(n2363)
  );


  SyncXor
  xor_C119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2363),
    .din1(n2364),
    .dout0(n2365)
  );


  SyncXor
  xor_C12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1359),
    .din0(n1360),
    .dout0(n1362)
  );


  SyncXor
  xor_C120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2385),
    .din0(n2386),
    .dout0(n2388)
  );


  SyncXor
  xor_C121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2387),
    .din0(n2388),
    .dout0(n2389)
  );


  SyncXor
  xor_C122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2399),
    .din1(n2400),
    .dout0(n2401)
  );


  SyncXor
  xor_C123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2401),
    .din1(n2402),
    .dout0(n2403)
  );


  SyncXor
  xor_C124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2423),
    .din0(n2424),
    .dout0(n2426)
  );


  SyncXor
  xor_C125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2425),
    .din0(n2426),
    .dout0(n2427)
  );


  SyncXor
  xor_C126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2437),
    .din1(n2438),
    .dout0(n2439)
  );


  SyncXor
  xor_C127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2439),
    .din1(n2440),
    .dout0(n2441)
  );


  SyncXor
  xor_C13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1361),
    .din0(n1362),
    .dout0(n1363)
  );


  SyncXor
  xor_C14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1373),
    .din1(n1374),
    .dout0(n1375)
  );


  SyncXor
  xor_C15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1375),
    .din1(n1376),
    .dout0(n1377)
  );


  SyncXor
  xor_C16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1397),
    .din0(n1398),
    .dout0(n1400)
  );


  SyncXor
  xor_C17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1399),
    .din0(n1400),
    .dout0(n1401)
  );


  SyncXor
  xor_C18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1411),
    .din1(n1412),
    .dout0(n1413)
  );


  SyncXor
  xor_C19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1413),
    .din1(n1414),
    .dout0(n1415)
  );


  SyncXor
  xor_C2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1261),
    .din1(n1262),
    .dout0(n1263)
  );


  SyncXor
  xor_C20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1435),
    .din0(n1436),
    .dout0(n1438)
  );


  SyncXor
  xor_C21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1437),
    .din0(n1438),
    .dout0(n1439)
  );


  SyncXor
  xor_C22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1449),
    .din1(n1450),
    .dout0(n1451)
  );


  SyncXor
  xor_C23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1451),
    .din1(n1452),
    .dout0(n1453)
  );


  SyncXor
  xor_C24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1473),
    .din0(n1474),
    .dout0(n1476)
  );


  SyncXor
  xor_C25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1475),
    .din0(n1476),
    .dout0(n1477)
  );


  SyncXor
  xor_C26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1487),
    .din1(n1488),
    .dout0(n1489)
  );


  SyncXor
  xor_C27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1489),
    .din1(n1490),
    .dout0(n1491)
  );


  SyncXor
  xor_C28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1511),
    .din0(n1512),
    .dout0(n1514)
  );


  SyncXor
  xor_C29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1513),
    .din0(n1514),
    .dout0(n1515)
  );


  SyncXor
  xor_C3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1263),
    .din1(n1264),
    .dout0(n1265)
  );


  SyncXor
  xor_C30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1525),
    .din1(n1526),
    .dout0(n1527)
  );


  SyncXor
  xor_C31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1527),
    .din1(n1528),
    .dout0(n1529)
  );


  SyncXor
  xor_C32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1549),
    .din0(n1550),
    .dout0(n1552)
  );


  SyncXor
  xor_C33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1551),
    .din0(n1552),
    .dout0(n1553)
  );


  SyncXor
  xor_C34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1563),
    .din1(n1564),
    .dout0(n1565)
  );


  SyncXor
  xor_C35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1565),
    .din1(n1566),
    .dout0(n1567)
  );


  SyncXor
  xor_C36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1587),
    .din0(n1588),
    .dout0(n1590)
  );


  SyncXor
  xor_C37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1589),
    .din0(n1590),
    .dout0(n1591)
  );


  SyncXor
  xor_C38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1601),
    .din1(n1602),
    .dout0(n1603)
  );


  SyncXor
  xor_C39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1603),
    .din1(n1604),
    .dout0(n1605)
  );


  SyncXor
  xor_C4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1283),
    .din0(n1284),
    .dout0(n1286)
  );


  SyncXor
  xor_C40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1625),
    .din0(n1626),
    .dout0(n1628)
  );


  SyncXor
  xor_C41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1627),
    .din0(n1628),
    .dout0(n1629)
  );


  SyncXor
  xor_C42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1639),
    .din1(n1640),
    .dout0(n1641)
  );


  SyncXor
  xor_C43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1641),
    .din1(n1642),
    .dout0(n1643)
  );


  SyncXor
  xor_C44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1663),
    .din0(n1664),
    .dout0(n1666)
  );


  SyncXor
  xor_C45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1665),
    .din0(n1666),
    .dout0(n1667)
  );


  SyncXor
  xor_C46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1677),
    .din1(n1678),
    .dout0(n1679)
  );


  SyncXor
  xor_C47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1679),
    .din1(n1680),
    .dout0(n1681)
  );


  SyncXor
  xor_C48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1701),
    .din0(n1702),
    .dout0(n1704)
  );


  SyncXor
  xor_C49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1703),
    .din0(n1704),
    .dout0(n1705)
  );


  SyncXor
  xor_C5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1285),
    .din0(n1286),
    .dout0(n1287)
  );


  SyncXor
  xor_C50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1715),
    .din1(n1716),
    .dout0(n1717)
  );


  SyncXor
  xor_C51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1717),
    .din1(n1718),
    .dout0(n1719)
  );


  SyncXor
  xor_C52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1739),
    .din0(n1740),
    .dout0(n1742)
  );


  SyncXor
  xor_C53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1741),
    .din0(n1742),
    .dout0(n1743)
  );


  SyncXor
  xor_C54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1753),
    .din1(n1754),
    .dout0(n1755)
  );


  SyncXor
  xor_C55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1755),
    .din1(n1756),
    .dout0(n1757)
  );


  SyncXor
  xor_C56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1777),
    .din0(n1778),
    .dout0(n1780)
  );


  SyncXor
  xor_C57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1779),
    .din0(n1780),
    .dout0(n1781)
  );


  SyncXor
  xor_C58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1791),
    .din1(n1792),
    .dout0(n1793)
  );


  SyncXor
  xor_C59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1793),
    .din1(n1794),
    .dout0(n1795)
  );


  SyncXor
  xor_C6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1297),
    .din1(n1298),
    .dout0(n1299)
  );


  SyncXor
  xor_C60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1815),
    .din0(n1816),
    .dout0(n1818)
  );


  SyncXor
  xor_C61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1817),
    .din0(n1818),
    .dout0(n1819)
  );


  SyncXor
  xor_C62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1829),
    .din1(n1830),
    .dout0(n1831)
  );


  SyncXor
  xor_C63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1831),
    .din1(n1832),
    .dout0(n1833)
  );


  SyncXor
  xor_C64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1853),
    .din0(n1854),
    .dout0(n1856)
  );


  SyncXor
  xor_C65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1855),
    .din0(n1856),
    .dout0(n1857)
  );


  SyncXor
  xor_C66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1867),
    .din1(n1868),
    .dout0(n1869)
  );


  SyncXor
  xor_C67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1869),
    .din1(n1870),
    .dout0(n1871)
  );


  SyncXor
  xor_C68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1891),
    .din0(n1892),
    .dout0(n1894)
  );


  SyncXor
  xor_C69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1893),
    .din0(n1894),
    .dout0(n1895)
  );


  SyncXor
  xor_C7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1299),
    .din1(n1300),
    .dout0(n1301)
  );


  SyncXor
  xor_C70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1905),
    .din1(n1906),
    .dout0(n1907)
  );


  SyncXor
  xor_C71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1907),
    .din1(n1908),
    .dout0(n1909)
  );


  SyncXor
  xor_C72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1929),
    .din0(n1930),
    .dout0(n1932)
  );


  SyncXor
  xor_C73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1931),
    .din0(n1932),
    .dout0(n1933)
  );


  SyncXor
  xor_C74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1943),
    .din1(n1944),
    .dout0(n1945)
  );


  SyncXor
  xor_C75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1945),
    .din1(n1946),
    .dout0(n1947)
  );


  SyncXor
  xor_C76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1967),
    .din0(n1968),
    .dout0(n1970)
  );


  SyncXor
  xor_C77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1969),
    .din0(n1970),
    .dout0(n1971)
  );


  SyncXor
  xor_C78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1981),
    .din1(n1982),
    .dout0(n1983)
  );


  SyncXor
  xor_C79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1983),
    .din1(n1984),
    .dout0(n1985)
  );


  SyncXor
  xor_C8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1321),
    .din0(n1322),
    .dout0(n1324)
  );


  SyncXor
  xor_C80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2005),
    .din0(n2006),
    .dout0(n2008)
  );


  SyncXor
  xor_C81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2007),
    .din0(n2008),
    .dout0(n2009)
  );


  SyncXor
  xor_C82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2019),
    .din1(n2020),
    .dout0(n2021)
  );


  SyncXor
  xor_C83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2021),
    .din1(n2022),
    .dout0(n2023)
  );


  SyncXor
  xor_C84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2043),
    .din0(n2044),
    .dout0(n2046)
  );


  SyncXor
  xor_C85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2045),
    .din0(n2046),
    .dout0(n2047)
  );


  SyncXor
  xor_C86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2057),
    .din1(n2058),
    .dout0(n2059)
  );


  SyncXor
  xor_C87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2059),
    .din1(n2060),
    .dout0(n2061)
  );


  SyncXor
  xor_C88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2081),
    .din0(n2082),
    .dout0(n2084)
  );


  SyncXor
  xor_C89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2083),
    .din0(n2084),
    .dout0(n2085)
  );


  SyncXor
  xor_C9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1323),
    .din0(n1324),
    .dout0(n1325)
  );


  SyncXor
  xor_C90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2095),
    .din1(n2096),
    .dout0(n2097)
  );


  SyncXor
  xor_C91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2097),
    .din1(n2098),
    .dout0(n2099)
  );


  SyncXor
  xor_C92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2119),
    .din0(n2120),
    .dout0(n2122)
  );


  SyncXor
  xor_C93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2121),
    .din0(n2122),
    .dout0(n2123)
  );


  SyncXor
  xor_C94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2133),
    .din1(n2134),
    .dout0(n2135)
  );


  SyncXor
  xor_C95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2135),
    .din1(n2136),
    .dout0(n2137)
  );


  SyncXor
  xor_C96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2157),
    .din0(n2158),
    .dout0(n2160)
  );


  SyncXor
  xor_C97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n2159),
    .din0(n2160),
    .dout0(n2161)
  );


  SyncXor
  xor_C98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2171),
    .din1(n2172),
    .dout0(n2173)
  );


  SyncXor
  xor_C99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n2173),
    .din1(n2174),
    .dout0(n2175)
  );


  SyncXor
  xor_D0
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n17),
    .din0(n18),
    .dout0(n20)
  );


  SyncXor
  xor_D1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n19),
    .din0(n20),
    .dout0(n21)
  );


  SyncXor
  xor_D10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n105),
    .din1(n106),
    .dout0(n107)
  );


  SyncXor
  xor_D100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n965),
    .din0(n966),
    .dout0(n968)
  );


  SyncXor
  xor_D101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n967),
    .din0(n968),
    .dout0(n969)
  );


  SyncXor
  xor_D102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n979),
    .din1(n980),
    .dout0(n981)
  );


  SyncXor
  xor_D103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n981),
    .din1(n982),
    .dout0(n983)
  );


  SyncXor
  xor_D104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1003),
    .din0(n1004),
    .dout0(n1006)
  );


  SyncXor
  xor_D105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1005),
    .din0(n1006),
    .dout0(n1007)
  );


  SyncXor
  xor_D106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1017),
    .din1(n1018),
    .dout0(n1019)
  );


  SyncXor
  xor_D107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1019),
    .din1(n1020),
    .dout0(n1021)
  );


  SyncXor
  xor_D108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1041),
    .din0(n1042),
    .dout0(n1044)
  );


  SyncXor
  xor_D109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1043),
    .din0(n1044),
    .dout0(n1045)
  );


  SyncXor
  xor_D11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n107),
    .din1(n108),
    .dout0(n109)
  );


  SyncXor
  xor_D110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1055),
    .din1(n1056),
    .dout0(n1057)
  );


  SyncXor
  xor_D111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1057),
    .din1(n1058),
    .dout0(n1059)
  );


  SyncXor
  xor_D112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1079),
    .din0(n1080),
    .dout0(n1082)
  );


  SyncXor
  xor_D113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1081),
    .din0(n1082),
    .dout0(n1083)
  );


  SyncXor
  xor_D114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1093),
    .din1(n1094),
    .dout0(n1095)
  );


  SyncXor
  xor_D115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1095),
    .din1(n1096),
    .dout0(n1097)
  );


  SyncXor
  xor_D116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1117),
    .din0(n1118),
    .dout0(n1120)
  );


  SyncXor
  xor_D117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1119),
    .din0(n1120),
    .dout0(n1121)
  );


  SyncXor
  xor_D118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1131),
    .din1(n1132),
    .dout0(n1133)
  );


  SyncXor
  xor_D119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1133),
    .din1(n1134),
    .dout0(n1135)
  );


  SyncXor
  xor_D12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n129),
    .din0(n130),
    .dout0(n132)
  );


  SyncXor
  xor_D120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1155),
    .din0(n1156),
    .dout0(n1158)
  );


  SyncXor
  xor_D121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1157),
    .din0(n1158),
    .dout0(n1159)
  );


  SyncXor
  xor_D122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1169),
    .din1(n1170),
    .dout0(n1171)
  );


  SyncXor
  xor_D123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1171),
    .din1(n1172),
    .dout0(n1173)
  );


  SyncXor
  xor_D124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1193),
    .din0(n1194),
    .dout0(n1196)
  );


  SyncXor
  xor_D125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n1195),
    .din0(n1196),
    .dout0(n1197)
  );


  SyncXor
  xor_D126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1207),
    .din1(n1208),
    .dout0(n1209)
  );


  SyncXor
  xor_D127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n1209),
    .din1(n1210),
    .dout0(n1211)
  );


  SyncXor
  xor_D13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n131),
    .din0(n132),
    .dout0(n133)
  );


  SyncXor
  xor_D14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n143),
    .din1(n144),
    .dout0(n145)
  );


  SyncXor
  xor_D15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n145),
    .din1(n146),
    .dout0(n147)
  );


  SyncXor
  xor_D16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n167),
    .din0(n168),
    .dout0(n170)
  );


  SyncXor
  xor_D17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n169),
    .din0(n170),
    .dout0(n171)
  );


  SyncXor
  xor_D18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n181),
    .din1(n182),
    .dout0(n183)
  );


  SyncXor
  xor_D19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n183),
    .din1(n184),
    .dout0(n185)
  );


  SyncXor
  xor_D2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n31),
    .din1(n32),
    .dout0(n33)
  );


  SyncXor
  xor_D20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n205),
    .din0(n206),
    .dout0(n208)
  );


  SyncXor
  xor_D21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n207),
    .din0(n208),
    .dout0(n209)
  );


  SyncXor
  xor_D22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n219),
    .din1(n220),
    .dout0(n221)
  );


  SyncXor
  xor_D23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n221),
    .din1(n222),
    .dout0(n223)
  );


  SyncXor
  xor_D24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n243),
    .din0(n244),
    .dout0(n246)
  );


  SyncXor
  xor_D25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n245),
    .din0(n246),
    .dout0(n247)
  );


  SyncXor
  xor_D26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n257),
    .din1(n258),
    .dout0(n259)
  );


  SyncXor
  xor_D27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n259),
    .din1(n260),
    .dout0(n261)
  );


  SyncXor
  xor_D28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n281),
    .din0(n282),
    .dout0(n284)
  );


  SyncXor
  xor_D29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n283),
    .din0(n284),
    .dout0(n285)
  );


  SyncXor
  xor_D3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n33),
    .din1(n34),
    .dout0(n35)
  );


  SyncXor
  xor_D30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n295),
    .din1(n296),
    .dout0(n297)
  );


  SyncXor
  xor_D31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n297),
    .din1(n298),
    .dout0(n299)
  );


  SyncXor
  xor_D32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n319),
    .din0(n320),
    .dout0(n322)
  );


  SyncXor
  xor_D33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n321),
    .din0(n322),
    .dout0(n323)
  );


  SyncXor
  xor_D34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n333),
    .din1(n334),
    .dout0(n335)
  );


  SyncXor
  xor_D35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n335),
    .din1(n336),
    .dout0(n337)
  );


  SyncXor
  xor_D36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n357),
    .din0(n358),
    .dout0(n360)
  );


  SyncXor
  xor_D37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n359),
    .din0(n360),
    .dout0(n361)
  );


  SyncXor
  xor_D38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n371),
    .din1(n372),
    .dout0(n373)
  );


  SyncXor
  xor_D39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n373),
    .din1(n374),
    .dout0(n375)
  );


  SyncXor
  xor_D4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n53),
    .din0(n54),
    .dout0(n56)
  );


  SyncXor
  xor_D40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n395),
    .din0(n396),
    .dout0(n398)
  );


  SyncXor
  xor_D41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n397),
    .din0(n398),
    .dout0(n399)
  );


  SyncXor
  xor_D42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n409),
    .din1(n410),
    .dout0(n411)
  );


  SyncXor
  xor_D43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n411),
    .din1(n412),
    .dout0(n413)
  );


  SyncXor
  xor_D44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n433),
    .din0(n434),
    .dout0(n436)
  );


  SyncXor
  xor_D45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n435),
    .din0(n436),
    .dout0(n437)
  );


  SyncXor
  xor_D46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n447),
    .din1(n448),
    .dout0(n449)
  );


  SyncXor
  xor_D47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n449),
    .din1(n450),
    .dout0(n451)
  );


  SyncXor
  xor_D48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n471),
    .din0(n472),
    .dout0(n474)
  );


  SyncXor
  xor_D49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n473),
    .din0(n474),
    .dout0(n475)
  );


  SyncXor
  xor_D5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n55),
    .din0(n56),
    .dout0(n57)
  );


  SyncXor
  xor_D50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n485),
    .din1(n486),
    .dout0(n487)
  );


  SyncXor
  xor_D51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n487),
    .din1(n488),
    .dout0(n489)
  );


  SyncXor
  xor_D52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n509),
    .din0(n510),
    .dout0(n512)
  );


  SyncXor
  xor_D53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n511),
    .din0(n512),
    .dout0(n513)
  );


  SyncXor
  xor_D54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n523),
    .din1(n524),
    .dout0(n525)
  );


  SyncXor
  xor_D55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n525),
    .din1(n526),
    .dout0(n527)
  );


  SyncXor
  xor_D56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n547),
    .din0(n548),
    .dout0(n550)
  );


  SyncXor
  xor_D57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n549),
    .din0(n550),
    .dout0(n551)
  );


  SyncXor
  xor_D58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n561),
    .din1(n562),
    .dout0(n563)
  );


  SyncXor
  xor_D59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n563),
    .din1(n564),
    .dout0(n565)
  );


  SyncXor
  xor_D6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n67),
    .din1(n68),
    .dout0(n69)
  );


  SyncXor
  xor_D60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n585),
    .din0(n586),
    .dout0(n588)
  );


  SyncXor
  xor_D61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n587),
    .din0(n588),
    .dout0(n589)
  );


  SyncXor
  xor_D62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n599),
    .din1(n600),
    .dout0(n601)
  );


  SyncXor
  xor_D63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n601),
    .din1(n602),
    .dout0(n603)
  );


  SyncXor
  xor_D64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n623),
    .din0(n624),
    .dout0(n626)
  );


  SyncXor
  xor_D65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n625),
    .din0(n626),
    .dout0(n627)
  );


  SyncXor
  xor_D66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n637),
    .din1(n638),
    .dout0(n639)
  );


  SyncXor
  xor_D67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n639),
    .din1(n640),
    .dout0(n641)
  );


  SyncXor
  xor_D68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n661),
    .din0(n662),
    .dout0(n664)
  );


  SyncXor
  xor_D69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n663),
    .din0(n664),
    .dout0(n665)
  );


  SyncXor
  xor_D7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n69),
    .din1(n70),
    .dout0(n71)
  );


  SyncXor
  xor_D70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n675),
    .din1(n676),
    .dout0(n677)
  );


  SyncXor
  xor_D71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n677),
    .din1(n678),
    .dout0(n679)
  );


  SyncXor
  xor_D72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n699),
    .din0(n700),
    .dout0(n702)
  );


  SyncXor
  xor_D73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n701),
    .din0(n702),
    .dout0(n703)
  );


  SyncXor
  xor_D74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n713),
    .din1(n714),
    .dout0(n715)
  );


  SyncXor
  xor_D75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n715),
    .din1(n716),
    .dout0(n717)
  );


  SyncXor
  xor_D76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n737),
    .din0(n738),
    .dout0(n740)
  );


  SyncXor
  xor_D77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n739),
    .din0(n740),
    .dout0(n741)
  );


  SyncXor
  xor_D78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n751),
    .din1(n752),
    .dout0(n753)
  );


  SyncXor
  xor_D79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n753),
    .din1(n754),
    .dout0(n755)
  );


  SyncXor
  xor_D8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n91),
    .din0(n92),
    .dout0(n94)
  );


  SyncXor
  xor_D80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n775),
    .din0(n776),
    .dout0(n778)
  );


  SyncXor
  xor_D81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n777),
    .din0(n778),
    .dout0(n779)
  );


  SyncXor
  xor_D82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n789),
    .din1(n790),
    .dout0(n791)
  );


  SyncXor
  xor_D83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n791),
    .din1(n792),
    .dout0(n793)
  );


  SyncXor
  xor_D84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n813),
    .din0(n814),
    .dout0(n816)
  );


  SyncXor
  xor_D85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n815),
    .din0(n816),
    .dout0(n817)
  );


  SyncXor
  xor_D86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n827),
    .din1(n828),
    .dout0(n829)
  );


  SyncXor
  xor_D87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n829),
    .din1(n830),
    .dout0(n831)
  );


  SyncXor
  xor_D88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n851),
    .din0(n852),
    .dout0(n854)
  );


  SyncXor
  xor_D89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n853),
    .din0(n854),
    .dout0(n855)
  );


  SyncXor
  xor_D9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n93),
    .din0(n94),
    .dout0(n95)
  );


  SyncXor
  xor_D90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n865),
    .din1(n866),
    .dout0(n867)
  );


  SyncXor
  xor_D91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n867),
    .din1(n868),
    .dout0(n869)
  );


  SyncXor
  xor_D92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n889),
    .din0(n890),
    .dout0(n892)
  );


  SyncXor
  xor_D93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n891),
    .din0(n892),
    .dout0(n893)
  );


  SyncXor
  xor_D94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n903),
    .din1(n904),
    .dout0(n905)
  );


  SyncXor
  xor_D95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n905),
    .din1(n906),
    .dout0(n907)
  );


  SyncXor
  xor_D96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n927),
    .din0(n928),
    .dout0(n930)
  );


  SyncXor
  xor_D97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din1(n929),
    .din0(n930),
    .dout0(n931)
  );


  SyncXor
  xor_D98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n941),
    .din1(n942),
    .dout0(n943)
  );


  SyncXor
  xor_D99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .din0(n943),
    .din1(n944),
    .dout0(n945)
  );


endmodule
