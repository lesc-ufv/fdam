module reg_tree_4_66_2 #
(
  parameter DATA_WIDTH = 16
)
(
  input clk,
  input [DATA_WIDTH-1:0] in,
  output [DATA_WIDTH-1:0] out_0,
  output [DATA_WIDTH-1:0] out_1,
  output [DATA_WIDTH-1:0] out_2,
  output [DATA_WIDTH-1:0] out_3,
  output [DATA_WIDTH-1:0] out_4,
  output [DATA_WIDTH-1:0] out_5,
  output [DATA_WIDTH-1:0] out_6,
  output [DATA_WIDTH-1:0] out_7,
  output [DATA_WIDTH-1:0] out_8,
  output [DATA_WIDTH-1:0] out_9,
  output [DATA_WIDTH-1:0] out_10,
  output [DATA_WIDTH-1:0] out_11,
  output [DATA_WIDTH-1:0] out_12,
  output [DATA_WIDTH-1:0] out_13,
  output [DATA_WIDTH-1:0] out_14,
  output [DATA_WIDTH-1:0] out_15,
  output [DATA_WIDTH-1:0] out_16,
  output [DATA_WIDTH-1:0] out_17,
  output [DATA_WIDTH-1:0] out_18,
  output [DATA_WIDTH-1:0] out_19,
  output [DATA_WIDTH-1:0] out_20,
  output [DATA_WIDTH-1:0] out_21,
  output [DATA_WIDTH-1:0] out_22,
  output [DATA_WIDTH-1:0] out_23,
  output [DATA_WIDTH-1:0] out_24,
  output [DATA_WIDTH-1:0] out_25,
  output [DATA_WIDTH-1:0] out_26,
  output [DATA_WIDTH-1:0] out_27,
  output [DATA_WIDTH-1:0] out_28,
  output [DATA_WIDTH-1:0] out_29,
  output [DATA_WIDTH-1:0] out_30,
  output [DATA_WIDTH-1:0] out_31,
  output [DATA_WIDTH-1:0] out_32,
  output [DATA_WIDTH-1:0] out_33,
  output [DATA_WIDTH-1:0] out_34,
  output [DATA_WIDTH-1:0] out_35,
  output [DATA_WIDTH-1:0] out_36,
  output [DATA_WIDTH-1:0] out_37,
  output [DATA_WIDTH-1:0] out_38,
  output [DATA_WIDTH-1:0] out_39,
  output [DATA_WIDTH-1:0] out_40,
  output [DATA_WIDTH-1:0] out_41,
  output [DATA_WIDTH-1:0] out_42,
  output [DATA_WIDTH-1:0] out_43,
  output [DATA_WIDTH-1:0] out_44,
  output [DATA_WIDTH-1:0] out_45,
  output [DATA_WIDTH-1:0] out_46,
  output [DATA_WIDTH-1:0] out_47,
  output [DATA_WIDTH-1:0] out_48,
  output [DATA_WIDTH-1:0] out_49,
  output [DATA_WIDTH-1:0] out_50,
  output [DATA_WIDTH-1:0] out_51,
  output [DATA_WIDTH-1:0] out_52,
  output [DATA_WIDTH-1:0] out_53,
  output [DATA_WIDTH-1:0] out_54,
  output [DATA_WIDTH-1:0] out_55,
  output [DATA_WIDTH-1:0] out_56,
  output [DATA_WIDTH-1:0] out_57,
  output [DATA_WIDTH-1:0] out_58,
  output [DATA_WIDTH-1:0] out_59,
  output [DATA_WIDTH-1:0] out_60,
  output [DATA_WIDTH-1:0] out_61,
  output [DATA_WIDTH-1:0] out_62,
  output [DATA_WIDTH-1:0] out_63,
  output [DATA_WIDTH-1:0] out_64,
  output [DATA_WIDTH-1:0] out_65
);

  reg [DATA_WIDTH-1:0] r [0:223-1];
  integer i;

  initial begin
    for(i=0; i<223; i=i+1) begin
      r[i] = 0;
    end
  end



  always @(posedge clk) begin
    r[0] <= in;
    r[1] <= r[0];
    r[2] <= r[0];
    r[3] <= r[1];
    r[4] <= r[1];
    r[5] <= r[1];
    r[6] <= r[1];
    r[7] <= r[2];
    r[8] <= r[3];
    r[9] <= r[3];
    r[10] <= r[3];
    r[11] <= r[3];
    r[12] <= r[4];
    r[13] <= r[4];
    r[14] <= r[4];
    r[15] <= r[4];
    r[16] <= r[5];
    r[17] <= r[5];
    r[18] <= r[5];
    r[19] <= r[5];
    r[20] <= r[6];
    r[21] <= r[6];
    r[22] <= r[6];
    r[23] <= r[6];
    r[24] <= r[7];
    r[25] <= r[8];
    r[26] <= r[8];
    r[27] <= r[8];
    r[28] <= r[8];
    r[29] <= r[9];
    r[30] <= r[9];
    r[31] <= r[9];
    r[32] <= r[9];
    r[33] <= r[10];
    r[34] <= r[10];
    r[35] <= r[10];
    r[36] <= r[10];
    r[37] <= r[11];
    r[38] <= r[11];
    r[39] <= r[11];
    r[40] <= r[11];
    r[41] <= r[12];
    r[42] <= r[12];
    r[43] <= r[12];
    r[44] <= r[12];
    r[45] <= r[13];
    r[46] <= r[13];
    r[47] <= r[13];
    r[48] <= r[13];
    r[49] <= r[14];
    r[50] <= r[14];
    r[51] <= r[14];
    r[52] <= r[14];
    r[53] <= r[15];
    r[54] <= r[15];
    r[55] <= r[15];
    r[56] <= r[15];
    r[57] <= r[16];
    r[58] <= r[16];
    r[59] <= r[16];
    r[60] <= r[16];
    r[61] <= r[17];
    r[62] <= r[17];
    r[63] <= r[17];
    r[64] <= r[17];
    r[65] <= r[18];
    r[66] <= r[18];
    r[67] <= r[18];
    r[68] <= r[18];
    r[69] <= r[19];
    r[70] <= r[19];
    r[71] <= r[19];
    r[72] <= r[19];
    r[73] <= r[20];
    r[74] <= r[20];
    r[75] <= r[20];
    r[76] <= r[20];
    r[77] <= r[21];
    r[78] <= r[21];
    r[79] <= r[21];
    r[80] <= r[21];
    r[81] <= r[22];
    r[82] <= r[22];
    r[83] <= r[22];
    r[84] <= r[22];
    r[85] <= r[23];
    r[86] <= r[23];
    r[87] <= r[23];
    r[88] <= r[23];
    r[89] <= r[24];
    r[90] <= r[24];
    r[91] <= r[25];
    r[92] <= r[26];
    r[93] <= r[27];
    r[94] <= r[28];
    r[95] <= r[29];
    r[96] <= r[30];
    r[97] <= r[31];
    r[98] <= r[32];
    r[99] <= r[33];
    r[100] <= r[34];
    r[101] <= r[35];
    r[102] <= r[36];
    r[103] <= r[37];
    r[104] <= r[38];
    r[105] <= r[39];
    r[106] <= r[40];
    r[107] <= r[41];
    r[108] <= r[42];
    r[109] <= r[43];
    r[110] <= r[44];
    r[111] <= r[45];
    r[112] <= r[46];
    r[113] <= r[47];
    r[114] <= r[48];
    r[115] <= r[49];
    r[116] <= r[50];
    r[117] <= r[51];
    r[118] <= r[52];
    r[119] <= r[53];
    r[120] <= r[54];
    r[121] <= r[55];
    r[122] <= r[56];
    r[123] <= r[57];
    r[124] <= r[58];
    r[125] <= r[59];
    r[126] <= r[60];
    r[127] <= r[61];
    r[128] <= r[62];
    r[129] <= r[63];
    r[130] <= r[64];
    r[131] <= r[65];
    r[132] <= r[66];
    r[133] <= r[67];
    r[134] <= r[68];
    r[135] <= r[69];
    r[136] <= r[70];
    r[137] <= r[71];
    r[138] <= r[72];
    r[139] <= r[73];
    r[140] <= r[74];
    r[141] <= r[75];
    r[142] <= r[76];
    r[143] <= r[77];
    r[144] <= r[78];
    r[145] <= r[79];
    r[146] <= r[80];
    r[147] <= r[81];
    r[148] <= r[82];
    r[149] <= r[83];
    r[150] <= r[84];
    r[151] <= r[85];
    r[152] <= r[86];
    r[153] <= r[87];
    r[154] <= r[88];
    r[155] <= r[89];
    r[156] <= r[90];
    r[157] <= r[91];
    r[158] <= r[92];
    r[159] <= r[93];
    r[160] <= r[94];
    r[161] <= r[95];
    r[162] <= r[96];
    r[163] <= r[97];
    r[164] <= r[98];
    r[165] <= r[99];
    r[166] <= r[100];
    r[167] <= r[101];
    r[168] <= r[102];
    r[169] <= r[103];
    r[170] <= r[104];
    r[171] <= r[105];
    r[172] <= r[106];
    r[173] <= r[107];
    r[174] <= r[108];
    r[175] <= r[109];
    r[176] <= r[110];
    r[177] <= r[111];
    r[178] <= r[112];
    r[179] <= r[113];
    r[180] <= r[114];
    r[181] <= r[115];
    r[182] <= r[116];
    r[183] <= r[117];
    r[184] <= r[118];
    r[185] <= r[119];
    r[186] <= r[120];
    r[187] <= r[121];
    r[188] <= r[122];
    r[189] <= r[123];
    r[190] <= r[124];
    r[191] <= r[125];
    r[192] <= r[126];
    r[193] <= r[127];
    r[194] <= r[128];
    r[195] <= r[129];
    r[196] <= r[130];
    r[197] <= r[131];
    r[198] <= r[132];
    r[199] <= r[133];
    r[200] <= r[134];
    r[201] <= r[135];
    r[202] <= r[136];
    r[203] <= r[137];
    r[204] <= r[138];
    r[205] <= r[139];
    r[206] <= r[140];
    r[207] <= r[141];
    r[208] <= r[142];
    r[209] <= r[143];
    r[210] <= r[144];
    r[211] <= r[145];
    r[212] <= r[146];
    r[213] <= r[147];
    r[214] <= r[148];
    r[215] <= r[149];
    r[216] <= r[150];
    r[217] <= r[151];
    r[218] <= r[152];
    r[219] <= r[153];
    r[220] <= r[154];
    r[221] <= r[155];
    r[222] <= r[156];

  end

  assign out_0 = r[157];
  assign out_1 = r[158];
  assign out_2 = r[159];
  assign out_3 = r[160];
  assign out_4 = r[161];
  assign out_5 = r[162];
  assign out_6 = r[163];
  assign out_7 = r[164];
  assign out_8 = r[165];
  assign out_9 = r[166];
  assign out_10 = r[167];
  assign out_11 = r[168];
  assign out_12 = r[169];
  assign out_13 = r[170];
  assign out_14 = r[171];
  assign out_15 = r[172];
  assign out_16 = r[173];
  assign out_17 = r[174];
  assign out_18 = r[175];
  assign out_19 = r[176];
  assign out_20 = r[177];
  assign out_21 = r[178];
  assign out_22 = r[179];
  assign out_23 = r[180];
  assign out_24 = r[181];
  assign out_25 = r[182];
  assign out_26 = r[183];
  assign out_27 = r[184];
  assign out_28 = r[185];
  assign out_29 = r[186];
  assign out_30 = r[187];
  assign out_31 = r[188];
  assign out_32 = r[189];
  assign out_33 = r[190];
  assign out_34 = r[191];
  assign out_35 = r[192];
  assign out_36 = r[193];
  assign out_37 = r[194];
  assign out_38 = r[195];
  assign out_39 = r[196];
  assign out_40 = r[197];
  assign out_41 = r[198];
  assign out_42 = r[199];
  assign out_43 = r[200];
  assign out_44 = r[201];
  assign out_45 = r[202];
  assign out_46 = r[203];
  assign out_47 = r[204];
  assign out_48 = r[205];
  assign out_49 = r[206];
  assign out_50 = r[207];
  assign out_51 = r[208];
  assign out_52 = r[209];
  assign out_53 = r[210];
  assign out_54 = r[211];
  assign out_55 = r[212];
  assign out_56 = r[213];
  assign out_57 = r[214];
  assign out_58 = r[215];
  assign out_59 = r[216];
  assign out_60 = r[217];
  assign out_61 = r[218];
  assign out_62 = r[219];
  assign out_63 = r[220];
  assign out_64 = r[221];
  assign out_65 = r[222];

endmodule