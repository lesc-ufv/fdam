module cgra0_top
(
  input clk,
  input rst,
  input [128-1:0] pes_en,
  input [64-1:0] conf_bus_in,
  input [1280-1:0] net_en,
  input [256-1:0] en_pc_net,
  output [8-1:0] fifo_in_re,
  input [128-1:0] fifo_in_data,
  output [8-1:0] fifo_out_we,
  output [128-1:0] fifo_out_data
);


  wire [64-1:0] conf_bus_0;
  wire [64-1:0] conf_bus_1;
  wire [64-1:0] conf_bus_2;
  wire [64-1:0] conf_bus_3;
  wire [64-1:0] conf_bus_4;
  wire [64-1:0] conf_bus_5;
  wire [64-1:0] conf_bus_6;
  wire [64-1:0] conf_bus_7;
  wire [64-1:0] conf_bus_8;
  wire [64-1:0] conf_bus_9;
  wire [64-1:0] conf_bus_10;
  wire [64-1:0] conf_bus_11;
  wire [64-1:0] conf_bus_12;
  wire [64-1:0] conf_bus_13;
  wire [64-1:0] conf_bus_14;
  wire [64-1:0] conf_bus_15;
  wire [64-1:0] conf_bus_16;
  wire [64-1:0] conf_bus_17;
  wire [64-1:0] conf_bus_18;
  wire [64-1:0] conf_bus_19;
  wire [64-1:0] conf_bus_20;
  wire [64-1:0] conf_bus_21;
  wire [64-1:0] conf_bus_22;
  wire [64-1:0] conf_bus_23;
  wire [64-1:0] conf_bus_24;
  wire [64-1:0] conf_bus_25;
  wire [64-1:0] conf_bus_26;
  wire [64-1:0] conf_bus_27;
  wire [64-1:0] conf_bus_28;
  wire [64-1:0] conf_bus_29;
  wire [64-1:0] conf_bus_30;
  wire [64-1:0] conf_bus_31;
  wire [64-1:0] conf_bus_32;
  wire [64-1:0] conf_bus_33;
  wire [64-1:0] conf_bus_34;
  wire [64-1:0] conf_bus_35;
  wire [64-1:0] conf_bus_36;
  wire [64-1:0] conf_bus_37;
  wire [64-1:0] conf_bus_38;
  wire [64-1:0] conf_bus_39;
  wire [64-1:0] conf_bus_40;
  wire [64-1:0] conf_bus_41;
  wire [64-1:0] conf_bus_42;
  wire [64-1:0] conf_bus_43;
  wire [64-1:0] conf_bus_44;
  wire [64-1:0] conf_bus_45;
  wire [64-1:0] conf_bus_46;
  wire [64-1:0] conf_bus_47;
  wire [64-1:0] conf_bus_48;
  wire [64-1:0] conf_bus_49;
  wire [64-1:0] conf_bus_50;
  wire [64-1:0] conf_bus_51;
  wire [64-1:0] conf_bus_52;
  wire [64-1:0] conf_bus_53;
  wire [64-1:0] conf_bus_54;
  wire [64-1:0] conf_bus_55;
  wire [64-1:0] conf_bus_56;
  wire [64-1:0] conf_bus_57;
  wire [64-1:0] conf_bus_58;
  wire [64-1:0] conf_bus_59;
  wire [64-1:0] conf_bus_60;
  wire [64-1:0] conf_bus_61;
  wire [64-1:0] conf_bus_62;
  wire [64-1:0] conf_bus_63;
  wire [64-1:0] conf_bus_64;
  wire [64-1:0] conf_bus_65;
  wire [64-1:0] conf_bus_66;
  wire [64-1:0] conf_bus_67;
  wire [64-1:0] conf_bus_68;
  wire [64-1:0] conf_bus_69;
  wire [64-1:0] conf_bus_70;
  wire [64-1:0] conf_bus_71;
  wire [64-1:0] conf_bus_72;
  wire [64-1:0] conf_bus_73;
  wire [64-1:0] conf_bus_74;
  wire [64-1:0] conf_bus_75;
  wire [64-1:0] conf_bus_76;
  wire [64-1:0] conf_bus_77;
  wire [64-1:0] conf_bus_78;
  wire [64-1:0] conf_bus_79;
  wire [64-1:0] conf_bus_80;
  wire [64-1:0] conf_bus_81;
  wire [64-1:0] conf_bus_82;
  wire [64-1:0] conf_bus_83;
  wire [64-1:0] conf_bus_84;
  wire [64-1:0] conf_bus_85;
  wire [64-1:0] conf_bus_86;
  wire [64-1:0] conf_bus_87;
  wire [64-1:0] conf_bus_88;
  wire [64-1:0] conf_bus_89;
  wire [64-1:0] conf_bus_90;
  wire [64-1:0] conf_bus_91;
  wire [64-1:0] conf_bus_92;
  wire [64-1:0] conf_bus_93;
  wire [64-1:0] conf_bus_94;
  wire [64-1:0] conf_bus_95;
  wire [64-1:0] conf_bus_96;
  wire [64-1:0] conf_bus_97;
  wire [64-1:0] conf_bus_98;
  wire [64-1:0] conf_bus_99;
  wire [64-1:0] conf_bus_100;
  wire [64-1:0] conf_bus_101;
  wire [64-1:0] conf_bus_102;
  wire [64-1:0] conf_bus_103;
  wire [64-1:0] conf_bus_104;
  wire [64-1:0] conf_bus_105;
  wire [64-1:0] conf_bus_106;
  wire [64-1:0] conf_bus_107;
  wire [64-1:0] conf_bus_108;
  wire [64-1:0] conf_bus_109;
  wire [64-1:0] conf_bus_110;
  wire [64-1:0] conf_bus_111;
  wire [64-1:0] conf_bus_112;
  wire [64-1:0] conf_bus_113;
  wire [64-1:0] conf_bus_114;
  wire [64-1:0] conf_bus_115;
  wire [64-1:0] conf_bus_116;
  wire [64-1:0] conf_bus_117;
  wire [64-1:0] conf_bus_118;
  wire [64-1:0] conf_bus_119;
  wire [64-1:0] conf_bus_120;
  wire [64-1:0] conf_bus_121;
  wire [64-1:0] conf_bus_122;
  wire [64-1:0] conf_bus_123;
  wire [64-1:0] conf_bus_124;
  wire [64-1:0] conf_bus_125;
  wire [64-1:0] conf_bus_126;
  wire [64-1:0] conf_bus_127;
  wire [64-1:0] conf_bus_128;
  wire [64-1:0] conf_bus_129;
  wire [16-1:0] pe2neta_0;
  wire [16-1:0] pe2neta_1;
  wire [16-1:0] pe2neta_2;
  wire [16-1:0] pe2neta_3;
  wire [16-1:0] pe2neta_4;
  wire [16-1:0] pe2neta_5;
  wire [16-1:0] pe2neta_6;
  wire [16-1:0] pe2neta_7;
  wire [16-1:0] pe2neta_8;
  wire [16-1:0] pe2neta_9;
  wire [16-1:0] pe2neta_10;
  wire [16-1:0] pe2neta_11;
  wire [16-1:0] pe2neta_12;
  wire [16-1:0] pe2neta_13;
  wire [16-1:0] pe2neta_14;
  wire [16-1:0] pe2neta_15;
  wire [16-1:0] pe2neta_16;
  wire [16-1:0] pe2neta_17;
  wire [16-1:0] pe2neta_18;
  wire [16-1:0] pe2neta_19;
  wire [16-1:0] pe2neta_20;
  wire [16-1:0] pe2neta_21;
  wire [16-1:0] pe2neta_22;
  wire [16-1:0] pe2neta_23;
  wire [16-1:0] pe2neta_24;
  wire [16-1:0] pe2neta_25;
  wire [16-1:0] pe2neta_26;
  wire [16-1:0] pe2neta_27;
  wire [16-1:0] pe2neta_28;
  wire [16-1:0] pe2neta_29;
  wire [16-1:0] pe2neta_30;
  wire [16-1:0] pe2neta_31;
  wire [16-1:0] pe2neta_32;
  wire [16-1:0] pe2neta_33;
  wire [16-1:0] pe2neta_34;
  wire [16-1:0] pe2neta_35;
  wire [16-1:0] pe2neta_36;
  wire [16-1:0] pe2neta_37;
  wire [16-1:0] pe2neta_38;
  wire [16-1:0] pe2neta_39;
  wire [16-1:0] pe2neta_40;
  wire [16-1:0] pe2neta_41;
  wire [16-1:0] pe2neta_42;
  wire [16-1:0] pe2neta_43;
  wire [16-1:0] pe2neta_44;
  wire [16-1:0] pe2neta_45;
  wire [16-1:0] pe2neta_46;
  wire [16-1:0] pe2neta_47;
  wire [16-1:0] pe2neta_48;
  wire [16-1:0] pe2neta_49;
  wire [16-1:0] pe2neta_50;
  wire [16-1:0] pe2neta_51;
  wire [16-1:0] pe2neta_52;
  wire [16-1:0] pe2neta_53;
  wire [16-1:0] pe2neta_54;
  wire [16-1:0] pe2neta_55;
  wire [16-1:0] pe2neta_56;
  wire [16-1:0] pe2neta_57;
  wire [16-1:0] pe2neta_58;
  wire [16-1:0] pe2neta_59;
  wire [16-1:0] pe2neta_60;
  wire [16-1:0] pe2neta_61;
  wire [16-1:0] pe2neta_62;
  wire [16-1:0] pe2neta_63;
  wire [16-1:0] pe2neta_64;
  wire [16-1:0] pe2neta_65;
  wire [16-1:0] pe2neta_66;
  wire [16-1:0] pe2neta_67;
  wire [16-1:0] pe2neta_68;
  wire [16-1:0] pe2neta_69;
  wire [16-1:0] pe2neta_70;
  wire [16-1:0] pe2neta_71;
  wire [16-1:0] pe2neta_72;
  wire [16-1:0] pe2neta_73;
  wire [16-1:0] pe2neta_74;
  wire [16-1:0] pe2neta_75;
  wire [16-1:0] pe2neta_76;
  wire [16-1:0] pe2neta_77;
  wire [16-1:0] pe2neta_78;
  wire [16-1:0] pe2neta_79;
  wire [16-1:0] pe2neta_80;
  wire [16-1:0] pe2neta_81;
  wire [16-1:0] pe2neta_82;
  wire [16-1:0] pe2neta_83;
  wire [16-1:0] pe2neta_84;
  wire [16-1:0] pe2neta_85;
  wire [16-1:0] pe2neta_86;
  wire [16-1:0] pe2neta_87;
  wire [16-1:0] pe2neta_88;
  wire [16-1:0] pe2neta_89;
  wire [16-1:0] pe2neta_90;
  wire [16-1:0] pe2neta_91;
  wire [16-1:0] pe2neta_92;
  wire [16-1:0] pe2neta_93;
  wire [16-1:0] pe2neta_94;
  wire [16-1:0] pe2neta_95;
  wire [16-1:0] pe2neta_96;
  wire [16-1:0] pe2neta_97;
  wire [16-1:0] pe2neta_98;
  wire [16-1:0] pe2neta_99;
  wire [16-1:0] pe2neta_100;
  wire [16-1:0] pe2neta_101;
  wire [16-1:0] pe2neta_102;
  wire [16-1:0] pe2neta_103;
  wire [16-1:0] pe2neta_104;
  wire [16-1:0] pe2neta_105;
  wire [16-1:0] pe2neta_106;
  wire [16-1:0] pe2neta_107;
  wire [16-1:0] pe2neta_108;
  wire [16-1:0] pe2neta_109;
  wire [16-1:0] pe2neta_110;
  wire [16-1:0] pe2neta_111;
  wire [16-1:0] pe2neta_112;
  wire [16-1:0] pe2neta_113;
  wire [16-1:0] pe2neta_114;
  wire [16-1:0] pe2neta_115;
  wire [16-1:0] pe2neta_116;
  wire [16-1:0] pe2neta_117;
  wire [16-1:0] pe2neta_118;
  wire [16-1:0] pe2neta_119;
  wire [16-1:0] pe2neta_120;
  wire [16-1:0] pe2neta_121;
  wire [16-1:0] pe2neta_122;
  wire [16-1:0] pe2neta_123;
  wire [16-1:0] pe2neta_124;
  wire [16-1:0] pe2neta_125;
  wire [16-1:0] pe2neta_126;
  wire [16-1:0] pe2neta_127;
  wire [16-1:0] pe2netb_0;
  wire [16-1:0] pe2netb_1;
  wire [16-1:0] pe2netb_2;
  wire [16-1:0] pe2netb_3;
  wire [16-1:0] pe2netb_4;
  wire [16-1:0] pe2netb_5;
  wire [16-1:0] pe2netb_6;
  wire [16-1:0] pe2netb_7;
  wire [16-1:0] pe2netb_8;
  wire [16-1:0] pe2netb_9;
  wire [16-1:0] pe2netb_10;
  wire [16-1:0] pe2netb_11;
  wire [16-1:0] pe2netb_12;
  wire [16-1:0] pe2netb_13;
  wire [16-1:0] pe2netb_14;
  wire [16-1:0] pe2netb_15;
  wire [16-1:0] pe2netb_16;
  wire [16-1:0] pe2netb_17;
  wire [16-1:0] pe2netb_18;
  wire [16-1:0] pe2netb_19;
  wire [16-1:0] pe2netb_20;
  wire [16-1:0] pe2netb_21;
  wire [16-1:0] pe2netb_22;
  wire [16-1:0] pe2netb_23;
  wire [16-1:0] pe2netb_24;
  wire [16-1:0] pe2netb_25;
  wire [16-1:0] pe2netb_26;
  wire [16-1:0] pe2netb_27;
  wire [16-1:0] pe2netb_28;
  wire [16-1:0] pe2netb_29;
  wire [16-1:0] pe2netb_30;
  wire [16-1:0] pe2netb_31;
  wire [16-1:0] pe2netb_32;
  wire [16-1:0] pe2netb_33;
  wire [16-1:0] pe2netb_34;
  wire [16-1:0] pe2netb_35;
  wire [16-1:0] pe2netb_36;
  wire [16-1:0] pe2netb_37;
  wire [16-1:0] pe2netb_38;
  wire [16-1:0] pe2netb_39;
  wire [16-1:0] pe2netb_40;
  wire [16-1:0] pe2netb_41;
  wire [16-1:0] pe2netb_42;
  wire [16-1:0] pe2netb_43;
  wire [16-1:0] pe2netb_44;
  wire [16-1:0] pe2netb_45;
  wire [16-1:0] pe2netb_46;
  wire [16-1:0] pe2netb_47;
  wire [16-1:0] pe2netb_48;
  wire [16-1:0] pe2netb_49;
  wire [16-1:0] pe2netb_50;
  wire [16-1:0] pe2netb_51;
  wire [16-1:0] pe2netb_52;
  wire [16-1:0] pe2netb_53;
  wire [16-1:0] pe2netb_54;
  wire [16-1:0] pe2netb_55;
  wire [16-1:0] pe2netb_56;
  wire [16-1:0] pe2netb_57;
  wire [16-1:0] pe2netb_58;
  wire [16-1:0] pe2netb_59;
  wire [16-1:0] pe2netb_60;
  wire [16-1:0] pe2netb_61;
  wire [16-1:0] pe2netb_62;
  wire [16-1:0] pe2netb_63;
  wire [16-1:0] pe2netb_64;
  wire [16-1:0] pe2netb_65;
  wire [16-1:0] pe2netb_66;
  wire [16-1:0] pe2netb_67;
  wire [16-1:0] pe2netb_68;
  wire [16-1:0] pe2netb_69;
  wire [16-1:0] pe2netb_70;
  wire [16-1:0] pe2netb_71;
  wire [16-1:0] pe2netb_72;
  wire [16-1:0] pe2netb_73;
  wire [16-1:0] pe2netb_74;
  wire [16-1:0] pe2netb_75;
  wire [16-1:0] pe2netb_76;
  wire [16-1:0] pe2netb_77;
  wire [16-1:0] pe2netb_78;
  wire [16-1:0] pe2netb_79;
  wire [16-1:0] pe2netb_80;
  wire [16-1:0] pe2netb_81;
  wire [16-1:0] pe2netb_82;
  wire [16-1:0] pe2netb_83;
  wire [16-1:0] pe2netb_84;
  wire [16-1:0] pe2netb_85;
  wire [16-1:0] pe2netb_86;
  wire [16-1:0] pe2netb_87;
  wire [16-1:0] pe2netb_88;
  wire [16-1:0] pe2netb_89;
  wire [16-1:0] pe2netb_90;
  wire [16-1:0] pe2netb_91;
  wire [16-1:0] pe2netb_92;
  wire [16-1:0] pe2netb_93;
  wire [16-1:0] pe2netb_94;
  wire [16-1:0] pe2netb_95;
  wire [16-1:0] pe2netb_96;
  wire [16-1:0] pe2netb_97;
  wire [16-1:0] pe2netb_98;
  wire [16-1:0] pe2netb_99;
  wire [16-1:0] pe2netb_100;
  wire [16-1:0] pe2netb_101;
  wire [16-1:0] pe2netb_102;
  wire [16-1:0] pe2netb_103;
  wire [16-1:0] pe2netb_104;
  wire [16-1:0] pe2netb_105;
  wire [16-1:0] pe2netb_106;
  wire [16-1:0] pe2netb_107;
  wire [16-1:0] pe2netb_108;
  wire [16-1:0] pe2netb_109;
  wire [16-1:0] pe2netb_110;
  wire [16-1:0] pe2netb_111;
  wire [16-1:0] pe2netb_112;
  wire [16-1:0] pe2netb_113;
  wire [16-1:0] pe2netb_114;
  wire [16-1:0] pe2netb_115;
  wire [16-1:0] pe2netb_116;
  wire [16-1:0] pe2netb_117;
  wire [16-1:0] pe2netb_118;
  wire [16-1:0] pe2netb_119;
  wire [16-1:0] pe2netb_120;
  wire [16-1:0] pe2netb_121;
  wire [16-1:0] pe2netb_122;
  wire [16-1:0] pe2netb_123;
  wire [16-1:0] pe2netb_124;
  wire [16-1:0] pe2netb_125;
  wire [16-1:0] pe2netb_126;
  wire [16-1:0] pe2netb_127;
  wire [16-1:0] net2pea_0;
  wire [16-1:0] net2pea_1;
  wire [16-1:0] net2pea_2;
  wire [16-1:0] net2pea_3;
  wire [16-1:0] net2pea_4;
  wire [16-1:0] net2pea_5;
  wire [16-1:0] net2pea_6;
  wire [16-1:0] net2pea_7;
  wire [16-1:0] net2pea_8;
  wire [16-1:0] net2pea_9;
  wire [16-1:0] net2pea_10;
  wire [16-1:0] net2pea_11;
  wire [16-1:0] net2pea_12;
  wire [16-1:0] net2pea_13;
  wire [16-1:0] net2pea_14;
  wire [16-1:0] net2pea_15;
  wire [16-1:0] net2pea_16;
  wire [16-1:0] net2pea_17;
  wire [16-1:0] net2pea_18;
  wire [16-1:0] net2pea_19;
  wire [16-1:0] net2pea_20;
  wire [16-1:0] net2pea_21;
  wire [16-1:0] net2pea_22;
  wire [16-1:0] net2pea_23;
  wire [16-1:0] net2pea_24;
  wire [16-1:0] net2pea_25;
  wire [16-1:0] net2pea_26;
  wire [16-1:0] net2pea_27;
  wire [16-1:0] net2pea_28;
  wire [16-1:0] net2pea_29;
  wire [16-1:0] net2pea_30;
  wire [16-1:0] net2pea_31;
  wire [16-1:0] net2pea_32;
  wire [16-1:0] net2pea_33;
  wire [16-1:0] net2pea_34;
  wire [16-1:0] net2pea_35;
  wire [16-1:0] net2pea_36;
  wire [16-1:0] net2pea_37;
  wire [16-1:0] net2pea_38;
  wire [16-1:0] net2pea_39;
  wire [16-1:0] net2pea_40;
  wire [16-1:0] net2pea_41;
  wire [16-1:0] net2pea_42;
  wire [16-1:0] net2pea_43;
  wire [16-1:0] net2pea_44;
  wire [16-1:0] net2pea_45;
  wire [16-1:0] net2pea_46;
  wire [16-1:0] net2pea_47;
  wire [16-1:0] net2pea_48;
  wire [16-1:0] net2pea_49;
  wire [16-1:0] net2pea_50;
  wire [16-1:0] net2pea_51;
  wire [16-1:0] net2pea_52;
  wire [16-1:0] net2pea_53;
  wire [16-1:0] net2pea_54;
  wire [16-1:0] net2pea_55;
  wire [16-1:0] net2pea_56;
  wire [16-1:0] net2pea_57;
  wire [16-1:0] net2pea_58;
  wire [16-1:0] net2pea_59;
  wire [16-1:0] net2pea_60;
  wire [16-1:0] net2pea_61;
  wire [16-1:0] net2pea_62;
  wire [16-1:0] net2pea_63;
  wire [16-1:0] net2pea_64;
  wire [16-1:0] net2pea_65;
  wire [16-1:0] net2pea_66;
  wire [16-1:0] net2pea_67;
  wire [16-1:0] net2pea_68;
  wire [16-1:0] net2pea_69;
  wire [16-1:0] net2pea_70;
  wire [16-1:0] net2pea_71;
  wire [16-1:0] net2pea_72;
  wire [16-1:0] net2pea_73;
  wire [16-1:0] net2pea_74;
  wire [16-1:0] net2pea_75;
  wire [16-1:0] net2pea_76;
  wire [16-1:0] net2pea_77;
  wire [16-1:0] net2pea_78;
  wire [16-1:0] net2pea_79;
  wire [16-1:0] net2pea_80;
  wire [16-1:0] net2pea_81;
  wire [16-1:0] net2pea_82;
  wire [16-1:0] net2pea_83;
  wire [16-1:0] net2pea_84;
  wire [16-1:0] net2pea_85;
  wire [16-1:0] net2pea_86;
  wire [16-1:0] net2pea_87;
  wire [16-1:0] net2pea_88;
  wire [16-1:0] net2pea_89;
  wire [16-1:0] net2pea_90;
  wire [16-1:0] net2pea_91;
  wire [16-1:0] net2pea_92;
  wire [16-1:0] net2pea_93;
  wire [16-1:0] net2pea_94;
  wire [16-1:0] net2pea_95;
  wire [16-1:0] net2pea_96;
  wire [16-1:0] net2pea_97;
  wire [16-1:0] net2pea_98;
  wire [16-1:0] net2pea_99;
  wire [16-1:0] net2pea_100;
  wire [16-1:0] net2pea_101;
  wire [16-1:0] net2pea_102;
  wire [16-1:0] net2pea_103;
  wire [16-1:0] net2pea_104;
  wire [16-1:0] net2pea_105;
  wire [16-1:0] net2pea_106;
  wire [16-1:0] net2pea_107;
  wire [16-1:0] net2pea_108;
  wire [16-1:0] net2pea_109;
  wire [16-1:0] net2pea_110;
  wire [16-1:0] net2pea_111;
  wire [16-1:0] net2pea_112;
  wire [16-1:0] net2pea_113;
  wire [16-1:0] net2pea_114;
  wire [16-1:0] net2pea_115;
  wire [16-1:0] net2pea_116;
  wire [16-1:0] net2pea_117;
  wire [16-1:0] net2pea_118;
  wire [16-1:0] net2pea_119;
  wire [16-1:0] net2pea_120;
  wire [16-1:0] net2pea_121;
  wire [16-1:0] net2pea_122;
  wire [16-1:0] net2pea_123;
  wire [16-1:0] net2pea_124;
  wire [16-1:0] net2pea_125;
  wire [16-1:0] net2pea_126;
  wire [16-1:0] net2pea_127;
  wire [16-1:0] net2peb_0;
  wire [16-1:0] net2peb_1;
  wire [16-1:0] net2peb_2;
  wire [16-1:0] net2peb_3;
  wire [16-1:0] net2peb_4;
  wire [16-1:0] net2peb_5;
  wire [16-1:0] net2peb_6;
  wire [16-1:0] net2peb_7;
  wire [16-1:0] net2peb_8;
  wire [16-1:0] net2peb_9;
  wire [16-1:0] net2peb_10;
  wire [16-1:0] net2peb_11;
  wire [16-1:0] net2peb_12;
  wire [16-1:0] net2peb_13;
  wire [16-1:0] net2peb_14;
  wire [16-1:0] net2peb_15;
  wire [16-1:0] net2peb_16;
  wire [16-1:0] net2peb_17;
  wire [16-1:0] net2peb_18;
  wire [16-1:0] net2peb_19;
  wire [16-1:0] net2peb_20;
  wire [16-1:0] net2peb_21;
  wire [16-1:0] net2peb_22;
  wire [16-1:0] net2peb_23;
  wire [16-1:0] net2peb_24;
  wire [16-1:0] net2peb_25;
  wire [16-1:0] net2peb_26;
  wire [16-1:0] net2peb_27;
  wire [16-1:0] net2peb_28;
  wire [16-1:0] net2peb_29;
  wire [16-1:0] net2peb_30;
  wire [16-1:0] net2peb_31;
  wire [16-1:0] net2peb_32;
  wire [16-1:0] net2peb_33;
  wire [16-1:0] net2peb_34;
  wire [16-1:0] net2peb_35;
  wire [16-1:0] net2peb_36;
  wire [16-1:0] net2peb_37;
  wire [16-1:0] net2peb_38;
  wire [16-1:0] net2peb_39;
  wire [16-1:0] net2peb_40;
  wire [16-1:0] net2peb_41;
  wire [16-1:0] net2peb_42;
  wire [16-1:0] net2peb_43;
  wire [16-1:0] net2peb_44;
  wire [16-1:0] net2peb_45;
  wire [16-1:0] net2peb_46;
  wire [16-1:0] net2peb_47;
  wire [16-1:0] net2peb_48;
  wire [16-1:0] net2peb_49;
  wire [16-1:0] net2peb_50;
  wire [16-1:0] net2peb_51;
  wire [16-1:0] net2peb_52;
  wire [16-1:0] net2peb_53;
  wire [16-1:0] net2peb_54;
  wire [16-1:0] net2peb_55;
  wire [16-1:0] net2peb_56;
  wire [16-1:0] net2peb_57;
  wire [16-1:0] net2peb_58;
  wire [16-1:0] net2peb_59;
  wire [16-1:0] net2peb_60;
  wire [16-1:0] net2peb_61;
  wire [16-1:0] net2peb_62;
  wire [16-1:0] net2peb_63;
  wire [16-1:0] net2peb_64;
  wire [16-1:0] net2peb_65;
  wire [16-1:0] net2peb_66;
  wire [16-1:0] net2peb_67;
  wire [16-1:0] net2peb_68;
  wire [16-1:0] net2peb_69;
  wire [16-1:0] net2peb_70;
  wire [16-1:0] net2peb_71;
  wire [16-1:0] net2peb_72;
  wire [16-1:0] net2peb_73;
  wire [16-1:0] net2peb_74;
  wire [16-1:0] net2peb_75;
  wire [16-1:0] net2peb_76;
  wire [16-1:0] net2peb_77;
  wire [16-1:0] net2peb_78;
  wire [16-1:0] net2peb_79;
  wire [16-1:0] net2peb_80;
  wire [16-1:0] net2peb_81;
  wire [16-1:0] net2peb_82;
  wire [16-1:0] net2peb_83;
  wire [16-1:0] net2peb_84;
  wire [16-1:0] net2peb_85;
  wire [16-1:0] net2peb_86;
  wire [16-1:0] net2peb_87;
  wire [16-1:0] net2peb_88;
  wire [16-1:0] net2peb_89;
  wire [16-1:0] net2peb_90;
  wire [16-1:0] net2peb_91;
  wire [16-1:0] net2peb_92;
  wire [16-1:0] net2peb_93;
  wire [16-1:0] net2peb_94;
  wire [16-1:0] net2peb_95;
  wire [16-1:0] net2peb_96;
  wire [16-1:0] net2peb_97;
  wire [16-1:0] net2peb_98;
  wire [16-1:0] net2peb_99;
  wire [16-1:0] net2peb_100;
  wire [16-1:0] net2peb_101;
  wire [16-1:0] net2peb_102;
  wire [16-1:0] net2peb_103;
  wire [16-1:0] net2peb_104;
  wire [16-1:0] net2peb_105;
  wire [16-1:0] net2peb_106;
  wire [16-1:0] net2peb_107;
  wire [16-1:0] net2peb_108;
  wire [16-1:0] net2peb_109;
  wire [16-1:0] net2peb_110;
  wire [16-1:0] net2peb_111;
  wire [16-1:0] net2peb_112;
  wire [16-1:0] net2peb_113;
  wire [16-1:0] net2peb_114;
  wire [16-1:0] net2peb_115;
  wire [16-1:0] net2peb_116;
  wire [16-1:0] net2peb_117;
  wire [16-1:0] net2peb_118;
  wire [16-1:0] net2peb_119;
  wire [16-1:0] net2peb_120;
  wire [16-1:0] net2peb_121;
  wire [16-1:0] net2peb_122;
  wire [16-1:0] net2peb_123;
  wire [16-1:0] net2peb_124;
  wire [16-1:0] net2peb_125;
  wire [16-1:0] net2peb_126;
  wire [16-1:0] net2peb_127;
  wire pe2net_branch_0;
  wire pe2net_branch_1;
  wire pe2net_branch_2;
  wire pe2net_branch_3;
  wire pe2net_branch_4;
  wire pe2net_branch_5;
  wire pe2net_branch_6;
  wire pe2net_branch_7;
  wire pe2net_branch_8;
  wire pe2net_branch_9;
  wire pe2net_branch_10;
  wire pe2net_branch_11;
  wire pe2net_branch_12;
  wire pe2net_branch_13;
  wire pe2net_branch_14;
  wire pe2net_branch_15;
  wire pe2net_branch_16;
  wire pe2net_branch_17;
  wire pe2net_branch_18;
  wire pe2net_branch_19;
  wire pe2net_branch_20;
  wire pe2net_branch_21;
  wire pe2net_branch_22;
  wire pe2net_branch_23;
  wire pe2net_branch_24;
  wire pe2net_branch_25;
  wire pe2net_branch_26;
  wire pe2net_branch_27;
  wire pe2net_branch_28;
  wire pe2net_branch_29;
  wire pe2net_branch_30;
  wire pe2net_branch_31;
  wire pe2net_branch_32;
  wire pe2net_branch_33;
  wire pe2net_branch_34;
  wire pe2net_branch_35;
  wire pe2net_branch_36;
  wire pe2net_branch_37;
  wire pe2net_branch_38;
  wire pe2net_branch_39;
  wire pe2net_branch_40;
  wire pe2net_branch_41;
  wire pe2net_branch_42;
  wire pe2net_branch_43;
  wire pe2net_branch_44;
  wire pe2net_branch_45;
  wire pe2net_branch_46;
  wire pe2net_branch_47;
  wire pe2net_branch_48;
  wire pe2net_branch_49;
  wire pe2net_branch_50;
  wire pe2net_branch_51;
  wire pe2net_branch_52;
  wire pe2net_branch_53;
  wire pe2net_branch_54;
  wire pe2net_branch_55;
  wire pe2net_branch_56;
  wire pe2net_branch_57;
  wire pe2net_branch_58;
  wire pe2net_branch_59;
  wire pe2net_branch_60;
  wire pe2net_branch_61;
  wire pe2net_branch_62;
  wire pe2net_branch_63;
  wire pe2net_branch_64;
  wire pe2net_branch_65;
  wire pe2net_branch_66;
  wire pe2net_branch_67;
  wire pe2net_branch_68;
  wire pe2net_branch_69;
  wire pe2net_branch_70;
  wire pe2net_branch_71;
  wire pe2net_branch_72;
  wire pe2net_branch_73;
  wire pe2net_branch_74;
  wire pe2net_branch_75;
  wire pe2net_branch_76;
  wire pe2net_branch_77;
  wire pe2net_branch_78;
  wire pe2net_branch_79;
  wire pe2net_branch_80;
  wire pe2net_branch_81;
  wire pe2net_branch_82;
  wire pe2net_branch_83;
  wire pe2net_branch_84;
  wire pe2net_branch_85;
  wire pe2net_branch_86;
  wire pe2net_branch_87;
  wire pe2net_branch_88;
  wire pe2net_branch_89;
  wire pe2net_branch_90;
  wire pe2net_branch_91;
  wire pe2net_branch_92;
  wire pe2net_branch_93;
  wire pe2net_branch_94;
  wire pe2net_branch_95;
  wire pe2net_branch_96;
  wire pe2net_branch_97;
  wire pe2net_branch_98;
  wire pe2net_branch_99;
  wire pe2net_branch_100;
  wire pe2net_branch_101;
  wire pe2net_branch_102;
  wire pe2net_branch_103;
  wire pe2net_branch_104;
  wire pe2net_branch_105;
  wire pe2net_branch_106;
  wire pe2net_branch_107;
  wire pe2net_branch_108;
  wire pe2net_branch_109;
  wire pe2net_branch_110;
  wire pe2net_branch_111;
  wire pe2net_branch_112;
  wire pe2net_branch_113;
  wire pe2net_branch_114;
  wire pe2net_branch_115;
  wire pe2net_branch_116;
  wire pe2net_branch_117;
  wire pe2net_branch_118;
  wire pe2net_branch_119;
  wire pe2net_branch_120;
  wire pe2net_branch_121;
  wire pe2net_branch_122;
  wire pe2net_branch_123;
  wire pe2net_branch_124;
  wire pe2net_branch_125;
  wire pe2net_branch_126;
  wire pe2net_branch_127;
  wire net_branch2peb_0;
  wire net_branch2peb_1;
  wire net_branch2peb_2;
  wire net_branch2peb_3;
  wire net_branch2peb_4;
  wire net_branch2peb_5;
  wire net_branch2peb_6;
  wire net_branch2peb_7;
  wire net_branch2peb_8;
  wire net_branch2peb_9;
  wire net_branch2peb_10;
  wire net_branch2peb_11;
  wire net_branch2peb_12;
  wire net_branch2peb_13;
  wire net_branch2peb_14;
  wire net_branch2peb_15;
  wire net_branch2peb_16;
  wire net_branch2peb_17;
  wire net_branch2peb_18;
  wire net_branch2peb_19;
  wire net_branch2peb_20;
  wire net_branch2peb_21;
  wire net_branch2peb_22;
  wire net_branch2peb_23;
  wire net_branch2peb_24;
  wire net_branch2peb_25;
  wire net_branch2peb_26;
  wire net_branch2peb_27;
  wire net_branch2peb_28;
  wire net_branch2peb_29;
  wire net_branch2peb_30;
  wire net_branch2peb_31;
  wire net_branch2peb_32;
  wire net_branch2peb_33;
  wire net_branch2peb_34;
  wire net_branch2peb_35;
  wire net_branch2peb_36;
  wire net_branch2peb_37;
  wire net_branch2peb_38;
  wire net_branch2peb_39;
  wire net_branch2peb_40;
  wire net_branch2peb_41;
  wire net_branch2peb_42;
  wire net_branch2peb_43;
  wire net_branch2peb_44;
  wire net_branch2peb_45;
  wire net_branch2peb_46;
  wire net_branch2peb_47;
  wire net_branch2peb_48;
  wire net_branch2peb_49;
  wire net_branch2peb_50;
  wire net_branch2peb_51;
  wire net_branch2peb_52;
  wire net_branch2peb_53;
  wire net_branch2peb_54;
  wire net_branch2peb_55;
  wire net_branch2peb_56;
  wire net_branch2peb_57;
  wire net_branch2peb_58;
  wire net_branch2peb_59;
  wire net_branch2peb_60;
  wire net_branch2peb_61;
  wire net_branch2peb_62;
  wire net_branch2peb_63;
  wire net_branch2peb_64;
  wire net_branch2peb_65;
  wire net_branch2peb_66;
  wire net_branch2peb_67;
  wire net_branch2peb_68;
  wire net_branch2peb_69;
  wire net_branch2peb_70;
  wire net_branch2peb_71;
  wire net_branch2peb_72;
  wire net_branch2peb_73;
  wire net_branch2peb_74;
  wire net_branch2peb_75;
  wire net_branch2peb_76;
  wire net_branch2peb_77;
  wire net_branch2peb_78;
  wire net_branch2peb_79;
  wire net_branch2peb_80;
  wire net_branch2peb_81;
  wire net_branch2peb_82;
  wire net_branch2peb_83;
  wire net_branch2peb_84;
  wire net_branch2peb_85;
  wire net_branch2peb_86;
  wire net_branch2peb_87;
  wire net_branch2peb_88;
  wire net_branch2peb_89;
  wire net_branch2peb_90;
  wire net_branch2peb_91;
  wire net_branch2peb_92;
  wire net_branch2peb_93;
  wire net_branch2peb_94;
  wire net_branch2peb_95;
  wire net_branch2peb_96;
  wire net_branch2peb_97;
  wire net_branch2peb_98;
  wire net_branch2peb_99;
  wire net_branch2peb_100;
  wire net_branch2peb_101;
  wire net_branch2peb_102;
  wire net_branch2peb_103;
  wire net_branch2peb_104;
  wire net_branch2peb_105;
  wire net_branch2peb_106;
  wire net_branch2peb_107;
  wire net_branch2peb_108;
  wire net_branch2peb_109;
  wire net_branch2peb_110;
  wire net_branch2peb_111;
  wire net_branch2peb_112;
  wire net_branch2peb_113;
  wire net_branch2peb_114;
  wire net_branch2peb_115;
  wire net_branch2peb_116;
  wire net_branch2peb_117;
  wire net_branch2peb_118;
  wire net_branch2peb_119;
  wire net_branch2peb_120;
  wire net_branch2peb_121;
  wire net_branch2peb_122;
  wire net_branch2peb_123;
  wire net_branch2peb_124;
  wire net_branch2peb_125;
  wire net_branch2peb_126;
  wire net_branch2peb_127;


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  reg_conf_bus_in2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_in),
    .out(conf_bus_0)
  );


  cgra0_pe_in
  #(
    .PE_ID(1)
  )
  pe_io_in_1
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[0]),
    .conf_bus_in(conf_bus_0),
    .branch_in(net_branch2peb_0),
    .branch_out(pe2net_branch_0),
    .fifo_re(fifo_in_re[0]),
    .fifo_data(fifo_in_data[15:0]),
    .ina(net2pea_0),
    .inb(net2peb_0),
    .outa(pe2neta_0),
    .outb(pe2netb_0)
  );


  cgra0_pe_in
  #(
    .PE_ID(2)
  )
  pe_io_in_2
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[1]),
    .conf_bus_in(conf_bus_1),
    .branch_in(net_branch2peb_1),
    .branch_out(pe2net_branch_1),
    .fifo_re(fifo_in_re[1]),
    .fifo_data(fifo_in_data[31:16]),
    .ina(net2pea_1),
    .inb(net2peb_1),
    .outa(pe2neta_1),
    .outb(pe2netb_1)
  );


  cgra0_pe_in
  #(
    .PE_ID(3)
  )
  pe_io_in_3
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[2]),
    .conf_bus_in(conf_bus_2),
    .branch_in(net_branch2peb_2),
    .branch_out(pe2net_branch_2),
    .fifo_re(fifo_in_re[2]),
    .fifo_data(fifo_in_data[47:32]),
    .ina(net2pea_2),
    .inb(net2peb_2),
    .outa(pe2neta_2),
    .outb(pe2netb_2)
  );


  cgra0_pe_in
  #(
    .PE_ID(4)
  )
  pe_io_in_4
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[3]),
    .conf_bus_in(conf_bus_3),
    .branch_in(net_branch2peb_3),
    .branch_out(pe2net_branch_3),
    .fifo_re(fifo_in_re[3]),
    .fifo_data(fifo_in_data[63:48]),
    .ina(net2pea_3),
    .inb(net2peb_3),
    .outa(pe2neta_3),
    .outb(pe2netb_3)
  );


  cgra0_pe_in
  #(
    .PE_ID(5)
  )
  pe_io_in_5
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[4]),
    .conf_bus_in(conf_bus_4),
    .branch_in(net_branch2peb_4),
    .branch_out(pe2net_branch_4),
    .fifo_re(fifo_in_re[4]),
    .fifo_data(fifo_in_data[79:64]),
    .ina(net2pea_4),
    .inb(net2peb_4),
    .outa(pe2neta_4),
    .outb(pe2netb_4)
  );


  cgra0_pe_in
  #(
    .PE_ID(6)
  )
  pe_io_in_6
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[5]),
    .conf_bus_in(conf_bus_5),
    .branch_in(net_branch2peb_5),
    .branch_out(pe2net_branch_5),
    .fifo_re(fifo_in_re[5]),
    .fifo_data(fifo_in_data[95:80]),
    .ina(net2pea_5),
    .inb(net2peb_5),
    .outa(pe2neta_5),
    .outb(pe2netb_5)
  );


  cgra0_pe_in
  #(
    .PE_ID(7)
  )
  pe_io_in_7
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[6]),
    .conf_bus_in(conf_bus_6),
    .branch_in(net_branch2peb_6),
    .branch_out(pe2net_branch_6),
    .fifo_re(fifo_in_re[6]),
    .fifo_data(fifo_in_data[111:96]),
    .ina(net2pea_6),
    .inb(net2peb_6),
    .outa(pe2neta_6),
    .outb(pe2netb_6)
  );


  cgra0_pe_in
  #(
    .PE_ID(8)
  )
  pe_io_in_8
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[7]),
    .conf_bus_in(conf_bus_7),
    .branch_in(net_branch2peb_7),
    .branch_out(pe2net_branch_7),
    .fifo_re(fifo_in_re[7]),
    .fifo_data(fifo_in_data[127:112]),
    .ina(net2pea_7),
    .inb(net2peb_7),
    .outa(pe2neta_7),
    .outb(pe2netb_7)
  );


  cgra0_pe_out
  #(
    .PE_ID(9)
  )
  pe_io_out_9
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[8]),
    .conf_bus_in(conf_bus_8),
    .branch_in(net_branch2peb_8),
    .branch_out(pe2net_branch_8),
    .fifo_we(fifo_out_we[0]),
    .fifo_data(fifo_out_data[15:0]),
    .ina(net2pea_8),
    .inb(net2peb_8),
    .outa(pe2neta_8),
    .outb(pe2netb_8)
  );


  cgra0_pe_out
  #(
    .PE_ID(10)
  )
  pe_io_out_10
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[9]),
    .conf_bus_in(conf_bus_9),
    .branch_in(net_branch2peb_9),
    .branch_out(pe2net_branch_9),
    .fifo_we(fifo_out_we[1]),
    .fifo_data(fifo_out_data[31:16]),
    .ina(net2pea_9),
    .inb(net2peb_9),
    .outa(pe2neta_9),
    .outb(pe2netb_9)
  );


  cgra0_pe_out
  #(
    .PE_ID(11)
  )
  pe_io_out_11
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[10]),
    .conf_bus_in(conf_bus_10),
    .branch_in(net_branch2peb_10),
    .branch_out(pe2net_branch_10),
    .fifo_we(fifo_out_we[2]),
    .fifo_data(fifo_out_data[47:32]),
    .ina(net2pea_10),
    .inb(net2peb_10),
    .outa(pe2neta_10),
    .outb(pe2netb_10)
  );


  cgra0_pe_out
  #(
    .PE_ID(12)
  )
  pe_io_out_12
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[11]),
    .conf_bus_in(conf_bus_11),
    .branch_in(net_branch2peb_11),
    .branch_out(pe2net_branch_11),
    .fifo_we(fifo_out_we[3]),
    .fifo_data(fifo_out_data[63:48]),
    .ina(net2pea_11),
    .inb(net2peb_11),
    .outa(pe2neta_11),
    .outb(pe2netb_11)
  );


  cgra0_pe_out
  #(
    .PE_ID(13)
  )
  pe_io_out_13
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[12]),
    .conf_bus_in(conf_bus_12),
    .branch_in(net_branch2peb_12),
    .branch_out(pe2net_branch_12),
    .fifo_we(fifo_out_we[4]),
    .fifo_data(fifo_out_data[79:64]),
    .ina(net2pea_12),
    .inb(net2peb_12),
    .outa(pe2neta_12),
    .outb(pe2netb_12)
  );


  cgra0_pe_out
  #(
    .PE_ID(14)
  )
  pe_io_out_14
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[13]),
    .conf_bus_in(conf_bus_13),
    .branch_in(net_branch2peb_13),
    .branch_out(pe2net_branch_13),
    .fifo_we(fifo_out_we[5]),
    .fifo_data(fifo_out_data[95:80]),
    .ina(net2pea_13),
    .inb(net2peb_13),
    .outa(pe2neta_13),
    .outb(pe2netb_13)
  );


  cgra0_pe_out
  #(
    .PE_ID(15)
  )
  pe_io_out_15
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[14]),
    .conf_bus_in(conf_bus_14),
    .branch_in(net_branch2peb_14),
    .branch_out(pe2net_branch_14),
    .fifo_we(fifo_out_we[6]),
    .fifo_data(fifo_out_data[111:96]),
    .ina(net2pea_14),
    .inb(net2peb_14),
    .outa(pe2neta_14),
    .outb(pe2netb_14)
  );


  cgra0_pe_out
  #(
    .PE_ID(16)
  )
  pe_io_out_16
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[15]),
    .conf_bus_in(conf_bus_15),
    .branch_in(net_branch2peb_15),
    .branch_out(pe2net_branch_15),
    .fifo_we(fifo_out_we[7]),
    .fifo_data(fifo_out_data[127:112]),
    .ina(net2pea_15),
    .inb(net2peb_15),
    .outa(pe2neta_15),
    .outb(pe2netb_15)
  );


  cgra0_pe
  #(
    .PE_ID(17)
  )
  pe_17
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[16]),
    .conf_bus_in(conf_bus_16),
    .branch_in(net_branch2peb_16),
    .branch_out(pe2net_branch_16),
    .ina(net2pea_16),
    .inb(net2peb_16),
    .outa(pe2neta_16),
    .outb(pe2netb_16)
  );


  cgra0_pe
  #(
    .PE_ID(18)
  )
  pe_18
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[17]),
    .conf_bus_in(conf_bus_17),
    .branch_in(net_branch2peb_17),
    .branch_out(pe2net_branch_17),
    .ina(net2pea_17),
    .inb(net2peb_17),
    .outa(pe2neta_17),
    .outb(pe2netb_17)
  );


  cgra0_pe
  #(
    .PE_ID(19)
  )
  pe_19
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[18]),
    .conf_bus_in(conf_bus_18),
    .branch_in(net_branch2peb_18),
    .branch_out(pe2net_branch_18),
    .ina(net2pea_18),
    .inb(net2peb_18),
    .outa(pe2neta_18),
    .outb(pe2netb_18)
  );


  cgra0_pe
  #(
    .PE_ID(20)
  )
  pe_20
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[19]),
    .conf_bus_in(conf_bus_19),
    .branch_in(net_branch2peb_19),
    .branch_out(pe2net_branch_19),
    .ina(net2pea_19),
    .inb(net2peb_19),
    .outa(pe2neta_19),
    .outb(pe2netb_19)
  );


  cgra0_pe
  #(
    .PE_ID(21)
  )
  pe_21
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[20]),
    .conf_bus_in(conf_bus_20),
    .branch_in(net_branch2peb_20),
    .branch_out(pe2net_branch_20),
    .ina(net2pea_20),
    .inb(net2peb_20),
    .outa(pe2neta_20),
    .outb(pe2netb_20)
  );


  cgra0_pe
  #(
    .PE_ID(22)
  )
  pe_22
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[21]),
    .conf_bus_in(conf_bus_21),
    .branch_in(net_branch2peb_21),
    .branch_out(pe2net_branch_21),
    .ina(net2pea_21),
    .inb(net2peb_21),
    .outa(pe2neta_21),
    .outb(pe2netb_21)
  );


  cgra0_pe
  #(
    .PE_ID(23)
  )
  pe_23
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[22]),
    .conf_bus_in(conf_bus_22),
    .branch_in(net_branch2peb_22),
    .branch_out(pe2net_branch_22),
    .ina(net2pea_22),
    .inb(net2peb_22),
    .outa(pe2neta_22),
    .outb(pe2netb_22)
  );


  cgra0_pe
  #(
    .PE_ID(24)
  )
  pe_24
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[23]),
    .conf_bus_in(conf_bus_23),
    .branch_in(net_branch2peb_23),
    .branch_out(pe2net_branch_23),
    .ina(net2pea_23),
    .inb(net2peb_23),
    .outa(pe2neta_23),
    .outb(pe2netb_23)
  );


  cgra0_pe
  #(
    .PE_ID(25)
  )
  pe_25
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[24]),
    .conf_bus_in(conf_bus_24),
    .branch_in(net_branch2peb_24),
    .branch_out(pe2net_branch_24),
    .ina(net2pea_24),
    .inb(net2peb_24),
    .outa(pe2neta_24),
    .outb(pe2netb_24)
  );


  cgra0_pe
  #(
    .PE_ID(26)
  )
  pe_26
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[25]),
    .conf_bus_in(conf_bus_25),
    .branch_in(net_branch2peb_25),
    .branch_out(pe2net_branch_25),
    .ina(net2pea_25),
    .inb(net2peb_25),
    .outa(pe2neta_25),
    .outb(pe2netb_25)
  );


  cgra0_pe
  #(
    .PE_ID(27)
  )
  pe_27
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[26]),
    .conf_bus_in(conf_bus_26),
    .branch_in(net_branch2peb_26),
    .branch_out(pe2net_branch_26),
    .ina(net2pea_26),
    .inb(net2peb_26),
    .outa(pe2neta_26),
    .outb(pe2netb_26)
  );


  cgra0_pe
  #(
    .PE_ID(28)
  )
  pe_28
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[27]),
    .conf_bus_in(conf_bus_27),
    .branch_in(net_branch2peb_27),
    .branch_out(pe2net_branch_27),
    .ina(net2pea_27),
    .inb(net2peb_27),
    .outa(pe2neta_27),
    .outb(pe2netb_27)
  );


  cgra0_pe
  #(
    .PE_ID(29)
  )
  pe_29
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[28]),
    .conf_bus_in(conf_bus_28),
    .branch_in(net_branch2peb_28),
    .branch_out(pe2net_branch_28),
    .ina(net2pea_28),
    .inb(net2peb_28),
    .outa(pe2neta_28),
    .outb(pe2netb_28)
  );


  cgra0_pe
  #(
    .PE_ID(30)
  )
  pe_30
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[29]),
    .conf_bus_in(conf_bus_29),
    .branch_in(net_branch2peb_29),
    .branch_out(pe2net_branch_29),
    .ina(net2pea_29),
    .inb(net2peb_29),
    .outa(pe2neta_29),
    .outb(pe2netb_29)
  );


  cgra0_pe
  #(
    .PE_ID(31)
  )
  pe_31
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[30]),
    .conf_bus_in(conf_bus_30),
    .branch_in(net_branch2peb_30),
    .branch_out(pe2net_branch_30),
    .ina(net2pea_30),
    .inb(net2peb_30),
    .outa(pe2neta_30),
    .outb(pe2netb_30)
  );


  cgra0_pe
  #(
    .PE_ID(32)
  )
  pe_32
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[31]),
    .conf_bus_in(conf_bus_31),
    .branch_in(net_branch2peb_31),
    .branch_out(pe2net_branch_31),
    .ina(net2pea_31),
    .inb(net2peb_31),
    .outa(pe2neta_31),
    .outb(pe2netb_31)
  );


  cgra0_pe
  #(
    .PE_ID(33)
  )
  pe_33
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[32]),
    .conf_bus_in(conf_bus_32),
    .branch_in(net_branch2peb_32),
    .branch_out(pe2net_branch_32),
    .ina(net2pea_32),
    .inb(net2peb_32),
    .outa(pe2neta_32),
    .outb(pe2netb_32)
  );


  cgra0_pe
  #(
    .PE_ID(34)
  )
  pe_34
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[33]),
    .conf_bus_in(conf_bus_33),
    .branch_in(net_branch2peb_33),
    .branch_out(pe2net_branch_33),
    .ina(net2pea_33),
    .inb(net2peb_33),
    .outa(pe2neta_33),
    .outb(pe2netb_33)
  );


  cgra0_pe
  #(
    .PE_ID(35)
  )
  pe_35
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[34]),
    .conf_bus_in(conf_bus_34),
    .branch_in(net_branch2peb_34),
    .branch_out(pe2net_branch_34),
    .ina(net2pea_34),
    .inb(net2peb_34),
    .outa(pe2neta_34),
    .outb(pe2netb_34)
  );


  cgra0_pe
  #(
    .PE_ID(36)
  )
  pe_36
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[35]),
    .conf_bus_in(conf_bus_35),
    .branch_in(net_branch2peb_35),
    .branch_out(pe2net_branch_35),
    .ina(net2pea_35),
    .inb(net2peb_35),
    .outa(pe2neta_35),
    .outb(pe2netb_35)
  );


  cgra0_pe
  #(
    .PE_ID(37)
  )
  pe_37
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[36]),
    .conf_bus_in(conf_bus_36),
    .branch_in(net_branch2peb_36),
    .branch_out(pe2net_branch_36),
    .ina(net2pea_36),
    .inb(net2peb_36),
    .outa(pe2neta_36),
    .outb(pe2netb_36)
  );


  cgra0_pe
  #(
    .PE_ID(38)
  )
  pe_38
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[37]),
    .conf_bus_in(conf_bus_37),
    .branch_in(net_branch2peb_37),
    .branch_out(pe2net_branch_37),
    .ina(net2pea_37),
    .inb(net2peb_37),
    .outa(pe2neta_37),
    .outb(pe2netb_37)
  );


  cgra0_pe
  #(
    .PE_ID(39)
  )
  pe_39
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[38]),
    .conf_bus_in(conf_bus_38),
    .branch_in(net_branch2peb_38),
    .branch_out(pe2net_branch_38),
    .ina(net2pea_38),
    .inb(net2peb_38),
    .outa(pe2neta_38),
    .outb(pe2netb_38)
  );


  cgra0_pe
  #(
    .PE_ID(40)
  )
  pe_40
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[39]),
    .conf_bus_in(conf_bus_39),
    .branch_in(net_branch2peb_39),
    .branch_out(pe2net_branch_39),
    .ina(net2pea_39),
    .inb(net2peb_39),
    .outa(pe2neta_39),
    .outb(pe2netb_39)
  );


  cgra0_pe
  #(
    .PE_ID(41)
  )
  pe_41
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[40]),
    .conf_bus_in(conf_bus_40),
    .branch_in(net_branch2peb_40),
    .branch_out(pe2net_branch_40),
    .ina(net2pea_40),
    .inb(net2peb_40),
    .outa(pe2neta_40),
    .outb(pe2netb_40)
  );


  cgra0_pe
  #(
    .PE_ID(42)
  )
  pe_42
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[41]),
    .conf_bus_in(conf_bus_41),
    .branch_in(net_branch2peb_41),
    .branch_out(pe2net_branch_41),
    .ina(net2pea_41),
    .inb(net2peb_41),
    .outa(pe2neta_41),
    .outb(pe2netb_41)
  );


  cgra0_pe
  #(
    .PE_ID(43)
  )
  pe_43
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[42]),
    .conf_bus_in(conf_bus_42),
    .branch_in(net_branch2peb_42),
    .branch_out(pe2net_branch_42),
    .ina(net2pea_42),
    .inb(net2peb_42),
    .outa(pe2neta_42),
    .outb(pe2netb_42)
  );


  cgra0_pe
  #(
    .PE_ID(44)
  )
  pe_44
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[43]),
    .conf_bus_in(conf_bus_43),
    .branch_in(net_branch2peb_43),
    .branch_out(pe2net_branch_43),
    .ina(net2pea_43),
    .inb(net2peb_43),
    .outa(pe2neta_43),
    .outb(pe2netb_43)
  );


  cgra0_pe
  #(
    .PE_ID(45)
  )
  pe_45
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[44]),
    .conf_bus_in(conf_bus_44),
    .branch_in(net_branch2peb_44),
    .branch_out(pe2net_branch_44),
    .ina(net2pea_44),
    .inb(net2peb_44),
    .outa(pe2neta_44),
    .outb(pe2netb_44)
  );


  cgra0_pe
  #(
    .PE_ID(46)
  )
  pe_46
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[45]),
    .conf_bus_in(conf_bus_45),
    .branch_in(net_branch2peb_45),
    .branch_out(pe2net_branch_45),
    .ina(net2pea_45),
    .inb(net2peb_45),
    .outa(pe2neta_45),
    .outb(pe2netb_45)
  );


  cgra0_pe
  #(
    .PE_ID(47)
  )
  pe_47
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[46]),
    .conf_bus_in(conf_bus_46),
    .branch_in(net_branch2peb_46),
    .branch_out(pe2net_branch_46),
    .ina(net2pea_46),
    .inb(net2peb_46),
    .outa(pe2neta_46),
    .outb(pe2netb_46)
  );


  cgra0_pe
  #(
    .PE_ID(48)
  )
  pe_48
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[47]),
    .conf_bus_in(conf_bus_47),
    .branch_in(net_branch2peb_47),
    .branch_out(pe2net_branch_47),
    .ina(net2pea_47),
    .inb(net2peb_47),
    .outa(pe2neta_47),
    .outb(pe2netb_47)
  );


  cgra0_pe
  #(
    .PE_ID(49)
  )
  pe_49
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[48]),
    .conf_bus_in(conf_bus_48),
    .branch_in(net_branch2peb_48),
    .branch_out(pe2net_branch_48),
    .ina(net2pea_48),
    .inb(net2peb_48),
    .outa(pe2neta_48),
    .outb(pe2netb_48)
  );


  cgra0_pe
  #(
    .PE_ID(50)
  )
  pe_50
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[49]),
    .conf_bus_in(conf_bus_49),
    .branch_in(net_branch2peb_49),
    .branch_out(pe2net_branch_49),
    .ina(net2pea_49),
    .inb(net2peb_49),
    .outa(pe2neta_49),
    .outb(pe2netb_49)
  );


  cgra0_pe
  #(
    .PE_ID(51)
  )
  pe_51
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[50]),
    .conf_bus_in(conf_bus_50),
    .branch_in(net_branch2peb_50),
    .branch_out(pe2net_branch_50),
    .ina(net2pea_50),
    .inb(net2peb_50),
    .outa(pe2neta_50),
    .outb(pe2netb_50)
  );


  cgra0_pe
  #(
    .PE_ID(52)
  )
  pe_52
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[51]),
    .conf_bus_in(conf_bus_51),
    .branch_in(net_branch2peb_51),
    .branch_out(pe2net_branch_51),
    .ina(net2pea_51),
    .inb(net2peb_51),
    .outa(pe2neta_51),
    .outb(pe2netb_51)
  );


  cgra0_pe
  #(
    .PE_ID(53)
  )
  pe_53
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[52]),
    .conf_bus_in(conf_bus_52),
    .branch_in(net_branch2peb_52),
    .branch_out(pe2net_branch_52),
    .ina(net2pea_52),
    .inb(net2peb_52),
    .outa(pe2neta_52),
    .outb(pe2netb_52)
  );


  cgra0_pe
  #(
    .PE_ID(54)
  )
  pe_54
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[53]),
    .conf_bus_in(conf_bus_53),
    .branch_in(net_branch2peb_53),
    .branch_out(pe2net_branch_53),
    .ina(net2pea_53),
    .inb(net2peb_53),
    .outa(pe2neta_53),
    .outb(pe2netb_53)
  );


  cgra0_pe
  #(
    .PE_ID(55)
  )
  pe_55
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[54]),
    .conf_bus_in(conf_bus_54),
    .branch_in(net_branch2peb_54),
    .branch_out(pe2net_branch_54),
    .ina(net2pea_54),
    .inb(net2peb_54),
    .outa(pe2neta_54),
    .outb(pe2netb_54)
  );


  cgra0_pe
  #(
    .PE_ID(56)
  )
  pe_56
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[55]),
    .conf_bus_in(conf_bus_55),
    .branch_in(net_branch2peb_55),
    .branch_out(pe2net_branch_55),
    .ina(net2pea_55),
    .inb(net2peb_55),
    .outa(pe2neta_55),
    .outb(pe2netb_55)
  );


  cgra0_pe
  #(
    .PE_ID(57)
  )
  pe_57
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[56]),
    .conf_bus_in(conf_bus_56),
    .branch_in(net_branch2peb_56),
    .branch_out(pe2net_branch_56),
    .ina(net2pea_56),
    .inb(net2peb_56),
    .outa(pe2neta_56),
    .outb(pe2netb_56)
  );


  cgra0_pe
  #(
    .PE_ID(58)
  )
  pe_58
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[57]),
    .conf_bus_in(conf_bus_57),
    .branch_in(net_branch2peb_57),
    .branch_out(pe2net_branch_57),
    .ina(net2pea_57),
    .inb(net2peb_57),
    .outa(pe2neta_57),
    .outb(pe2netb_57)
  );


  cgra0_pe
  #(
    .PE_ID(59)
  )
  pe_59
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[58]),
    .conf_bus_in(conf_bus_58),
    .branch_in(net_branch2peb_58),
    .branch_out(pe2net_branch_58),
    .ina(net2pea_58),
    .inb(net2peb_58),
    .outa(pe2neta_58),
    .outb(pe2netb_58)
  );


  cgra0_pe
  #(
    .PE_ID(60)
  )
  pe_60
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[59]),
    .conf_bus_in(conf_bus_59),
    .branch_in(net_branch2peb_59),
    .branch_out(pe2net_branch_59),
    .ina(net2pea_59),
    .inb(net2peb_59),
    .outa(pe2neta_59),
    .outb(pe2netb_59)
  );


  cgra0_pe
  #(
    .PE_ID(61)
  )
  pe_61
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[60]),
    .conf_bus_in(conf_bus_60),
    .branch_in(net_branch2peb_60),
    .branch_out(pe2net_branch_60),
    .ina(net2pea_60),
    .inb(net2peb_60),
    .outa(pe2neta_60),
    .outb(pe2netb_60)
  );


  cgra0_pe
  #(
    .PE_ID(62)
  )
  pe_62
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[61]),
    .conf_bus_in(conf_bus_61),
    .branch_in(net_branch2peb_61),
    .branch_out(pe2net_branch_61),
    .ina(net2pea_61),
    .inb(net2peb_61),
    .outa(pe2neta_61),
    .outb(pe2netb_61)
  );


  cgra0_pe
  #(
    .PE_ID(63)
  )
  pe_63
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[62]),
    .conf_bus_in(conf_bus_62),
    .branch_in(net_branch2peb_62),
    .branch_out(pe2net_branch_62),
    .ina(net2pea_62),
    .inb(net2peb_62),
    .outa(pe2neta_62),
    .outb(pe2netb_62)
  );


  cgra0_pe
  #(
    .PE_ID(64)
  )
  pe_64
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[63]),
    .conf_bus_in(conf_bus_63),
    .branch_in(net_branch2peb_63),
    .branch_out(pe2net_branch_63),
    .ina(net2pea_63),
    .inb(net2peb_63),
    .outa(pe2neta_63),
    .outb(pe2netb_63)
  );


  cgra0_pe
  #(
    .PE_ID(65)
  )
  pe_65
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[64]),
    .conf_bus_in(conf_bus_64),
    .branch_in(net_branch2peb_64),
    .branch_out(pe2net_branch_64),
    .ina(net2pea_64),
    .inb(net2peb_64),
    .outa(pe2neta_64),
    .outb(pe2netb_64)
  );


  cgra0_pe
  #(
    .PE_ID(66)
  )
  pe_66
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[65]),
    .conf_bus_in(conf_bus_65),
    .branch_in(net_branch2peb_65),
    .branch_out(pe2net_branch_65),
    .ina(net2pea_65),
    .inb(net2peb_65),
    .outa(pe2neta_65),
    .outb(pe2netb_65)
  );


  cgra0_pe
  #(
    .PE_ID(67)
  )
  pe_67
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[66]),
    .conf_bus_in(conf_bus_66),
    .branch_in(net_branch2peb_66),
    .branch_out(pe2net_branch_66),
    .ina(net2pea_66),
    .inb(net2peb_66),
    .outa(pe2neta_66),
    .outb(pe2netb_66)
  );


  cgra0_pe
  #(
    .PE_ID(68)
  )
  pe_68
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[67]),
    .conf_bus_in(conf_bus_67),
    .branch_in(net_branch2peb_67),
    .branch_out(pe2net_branch_67),
    .ina(net2pea_67),
    .inb(net2peb_67),
    .outa(pe2neta_67),
    .outb(pe2netb_67)
  );


  cgra0_pe
  #(
    .PE_ID(69)
  )
  pe_69
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[68]),
    .conf_bus_in(conf_bus_68),
    .branch_in(net_branch2peb_68),
    .branch_out(pe2net_branch_68),
    .ina(net2pea_68),
    .inb(net2peb_68),
    .outa(pe2neta_68),
    .outb(pe2netb_68)
  );


  cgra0_pe
  #(
    .PE_ID(70)
  )
  pe_70
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[69]),
    .conf_bus_in(conf_bus_69),
    .branch_in(net_branch2peb_69),
    .branch_out(pe2net_branch_69),
    .ina(net2pea_69),
    .inb(net2peb_69),
    .outa(pe2neta_69),
    .outb(pe2netb_69)
  );


  cgra0_pe
  #(
    .PE_ID(71)
  )
  pe_71
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[70]),
    .conf_bus_in(conf_bus_70),
    .branch_in(net_branch2peb_70),
    .branch_out(pe2net_branch_70),
    .ina(net2pea_70),
    .inb(net2peb_70),
    .outa(pe2neta_70),
    .outb(pe2netb_70)
  );


  cgra0_pe
  #(
    .PE_ID(72)
  )
  pe_72
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[71]),
    .conf_bus_in(conf_bus_71),
    .branch_in(net_branch2peb_71),
    .branch_out(pe2net_branch_71),
    .ina(net2pea_71),
    .inb(net2peb_71),
    .outa(pe2neta_71),
    .outb(pe2netb_71)
  );


  cgra0_pe
  #(
    .PE_ID(73)
  )
  pe_73
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[72]),
    .conf_bus_in(conf_bus_72),
    .branch_in(net_branch2peb_72),
    .branch_out(pe2net_branch_72),
    .ina(net2pea_72),
    .inb(net2peb_72),
    .outa(pe2neta_72),
    .outb(pe2netb_72)
  );


  cgra0_pe
  #(
    .PE_ID(74)
  )
  pe_74
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[73]),
    .conf_bus_in(conf_bus_73),
    .branch_in(net_branch2peb_73),
    .branch_out(pe2net_branch_73),
    .ina(net2pea_73),
    .inb(net2peb_73),
    .outa(pe2neta_73),
    .outb(pe2netb_73)
  );


  cgra0_pe
  #(
    .PE_ID(75)
  )
  pe_75
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[74]),
    .conf_bus_in(conf_bus_74),
    .branch_in(net_branch2peb_74),
    .branch_out(pe2net_branch_74),
    .ina(net2pea_74),
    .inb(net2peb_74),
    .outa(pe2neta_74),
    .outb(pe2netb_74)
  );


  cgra0_pe
  #(
    .PE_ID(76)
  )
  pe_76
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[75]),
    .conf_bus_in(conf_bus_75),
    .branch_in(net_branch2peb_75),
    .branch_out(pe2net_branch_75),
    .ina(net2pea_75),
    .inb(net2peb_75),
    .outa(pe2neta_75),
    .outb(pe2netb_75)
  );


  cgra0_pe
  #(
    .PE_ID(77)
  )
  pe_77
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[76]),
    .conf_bus_in(conf_bus_76),
    .branch_in(net_branch2peb_76),
    .branch_out(pe2net_branch_76),
    .ina(net2pea_76),
    .inb(net2peb_76),
    .outa(pe2neta_76),
    .outb(pe2netb_76)
  );


  cgra0_pe
  #(
    .PE_ID(78)
  )
  pe_78
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[77]),
    .conf_bus_in(conf_bus_77),
    .branch_in(net_branch2peb_77),
    .branch_out(pe2net_branch_77),
    .ina(net2pea_77),
    .inb(net2peb_77),
    .outa(pe2neta_77),
    .outb(pe2netb_77)
  );


  cgra0_pe
  #(
    .PE_ID(79)
  )
  pe_79
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[78]),
    .conf_bus_in(conf_bus_78),
    .branch_in(net_branch2peb_78),
    .branch_out(pe2net_branch_78),
    .ina(net2pea_78),
    .inb(net2peb_78),
    .outa(pe2neta_78),
    .outb(pe2netb_78)
  );


  cgra0_pe
  #(
    .PE_ID(80)
  )
  pe_80
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[79]),
    .conf_bus_in(conf_bus_79),
    .branch_in(net_branch2peb_79),
    .branch_out(pe2net_branch_79),
    .ina(net2pea_79),
    .inb(net2peb_79),
    .outa(pe2neta_79),
    .outb(pe2netb_79)
  );


  cgra0_pe
  #(
    .PE_ID(81)
  )
  pe_81
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[80]),
    .conf_bus_in(conf_bus_80),
    .branch_in(net_branch2peb_80),
    .branch_out(pe2net_branch_80),
    .ina(net2pea_80),
    .inb(net2peb_80),
    .outa(pe2neta_80),
    .outb(pe2netb_80)
  );


  cgra0_pe
  #(
    .PE_ID(82)
  )
  pe_82
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[81]),
    .conf_bus_in(conf_bus_81),
    .branch_in(net_branch2peb_81),
    .branch_out(pe2net_branch_81),
    .ina(net2pea_81),
    .inb(net2peb_81),
    .outa(pe2neta_81),
    .outb(pe2netb_81)
  );


  cgra0_pe
  #(
    .PE_ID(83)
  )
  pe_83
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[82]),
    .conf_bus_in(conf_bus_82),
    .branch_in(net_branch2peb_82),
    .branch_out(pe2net_branch_82),
    .ina(net2pea_82),
    .inb(net2peb_82),
    .outa(pe2neta_82),
    .outb(pe2netb_82)
  );


  cgra0_pe
  #(
    .PE_ID(84)
  )
  pe_84
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[83]),
    .conf_bus_in(conf_bus_83),
    .branch_in(net_branch2peb_83),
    .branch_out(pe2net_branch_83),
    .ina(net2pea_83),
    .inb(net2peb_83),
    .outa(pe2neta_83),
    .outb(pe2netb_83)
  );


  cgra0_pe
  #(
    .PE_ID(85)
  )
  pe_85
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[84]),
    .conf_bus_in(conf_bus_84),
    .branch_in(net_branch2peb_84),
    .branch_out(pe2net_branch_84),
    .ina(net2pea_84),
    .inb(net2peb_84),
    .outa(pe2neta_84),
    .outb(pe2netb_84)
  );


  cgra0_pe
  #(
    .PE_ID(86)
  )
  pe_86
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[85]),
    .conf_bus_in(conf_bus_85),
    .branch_in(net_branch2peb_85),
    .branch_out(pe2net_branch_85),
    .ina(net2pea_85),
    .inb(net2peb_85),
    .outa(pe2neta_85),
    .outb(pe2netb_85)
  );


  cgra0_pe
  #(
    .PE_ID(87)
  )
  pe_87
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[86]),
    .conf_bus_in(conf_bus_86),
    .branch_in(net_branch2peb_86),
    .branch_out(pe2net_branch_86),
    .ina(net2pea_86),
    .inb(net2peb_86),
    .outa(pe2neta_86),
    .outb(pe2netb_86)
  );


  cgra0_pe
  #(
    .PE_ID(88)
  )
  pe_88
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[87]),
    .conf_bus_in(conf_bus_87),
    .branch_in(net_branch2peb_87),
    .branch_out(pe2net_branch_87),
    .ina(net2pea_87),
    .inb(net2peb_87),
    .outa(pe2neta_87),
    .outb(pe2netb_87)
  );


  cgra0_pe
  #(
    .PE_ID(89)
  )
  pe_89
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[88]),
    .conf_bus_in(conf_bus_88),
    .branch_in(net_branch2peb_88),
    .branch_out(pe2net_branch_88),
    .ina(net2pea_88),
    .inb(net2peb_88),
    .outa(pe2neta_88),
    .outb(pe2netb_88)
  );


  cgra0_pe
  #(
    .PE_ID(90)
  )
  pe_90
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[89]),
    .conf_bus_in(conf_bus_89),
    .branch_in(net_branch2peb_89),
    .branch_out(pe2net_branch_89),
    .ina(net2pea_89),
    .inb(net2peb_89),
    .outa(pe2neta_89),
    .outb(pe2netb_89)
  );


  cgra0_pe
  #(
    .PE_ID(91)
  )
  pe_91
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[90]),
    .conf_bus_in(conf_bus_90),
    .branch_in(net_branch2peb_90),
    .branch_out(pe2net_branch_90),
    .ina(net2pea_90),
    .inb(net2peb_90),
    .outa(pe2neta_90),
    .outb(pe2netb_90)
  );


  cgra0_pe
  #(
    .PE_ID(92)
  )
  pe_92
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[91]),
    .conf_bus_in(conf_bus_91),
    .branch_in(net_branch2peb_91),
    .branch_out(pe2net_branch_91),
    .ina(net2pea_91),
    .inb(net2peb_91),
    .outa(pe2neta_91),
    .outb(pe2netb_91)
  );


  cgra0_pe
  #(
    .PE_ID(93)
  )
  pe_93
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[92]),
    .conf_bus_in(conf_bus_92),
    .branch_in(net_branch2peb_92),
    .branch_out(pe2net_branch_92),
    .ina(net2pea_92),
    .inb(net2peb_92),
    .outa(pe2neta_92),
    .outb(pe2netb_92)
  );


  cgra0_pe
  #(
    .PE_ID(94)
  )
  pe_94
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[93]),
    .conf_bus_in(conf_bus_93),
    .branch_in(net_branch2peb_93),
    .branch_out(pe2net_branch_93),
    .ina(net2pea_93),
    .inb(net2peb_93),
    .outa(pe2neta_93),
    .outb(pe2netb_93)
  );


  cgra0_pe
  #(
    .PE_ID(95)
  )
  pe_95
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[94]),
    .conf_bus_in(conf_bus_94),
    .branch_in(net_branch2peb_94),
    .branch_out(pe2net_branch_94),
    .ina(net2pea_94),
    .inb(net2peb_94),
    .outa(pe2neta_94),
    .outb(pe2netb_94)
  );


  cgra0_pe
  #(
    .PE_ID(96)
  )
  pe_96
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[95]),
    .conf_bus_in(conf_bus_95),
    .branch_in(net_branch2peb_95),
    .branch_out(pe2net_branch_95),
    .ina(net2pea_95),
    .inb(net2peb_95),
    .outa(pe2neta_95),
    .outb(pe2netb_95)
  );


  cgra0_pe
  #(
    .PE_ID(97)
  )
  pe_97
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[96]),
    .conf_bus_in(conf_bus_96),
    .branch_in(net_branch2peb_96),
    .branch_out(pe2net_branch_96),
    .ina(net2pea_96),
    .inb(net2peb_96),
    .outa(pe2neta_96),
    .outb(pe2netb_96)
  );


  cgra0_pe
  #(
    .PE_ID(98)
  )
  pe_98
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[97]),
    .conf_bus_in(conf_bus_97),
    .branch_in(net_branch2peb_97),
    .branch_out(pe2net_branch_97),
    .ina(net2pea_97),
    .inb(net2peb_97),
    .outa(pe2neta_97),
    .outb(pe2netb_97)
  );


  cgra0_pe
  #(
    .PE_ID(99)
  )
  pe_99
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[98]),
    .conf_bus_in(conf_bus_98),
    .branch_in(net_branch2peb_98),
    .branch_out(pe2net_branch_98),
    .ina(net2pea_98),
    .inb(net2peb_98),
    .outa(pe2neta_98),
    .outb(pe2netb_98)
  );


  cgra0_pe
  #(
    .PE_ID(100)
  )
  pe_100
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[99]),
    .conf_bus_in(conf_bus_99),
    .branch_in(net_branch2peb_99),
    .branch_out(pe2net_branch_99),
    .ina(net2pea_99),
    .inb(net2peb_99),
    .outa(pe2neta_99),
    .outb(pe2netb_99)
  );


  cgra0_pe
  #(
    .PE_ID(101)
  )
  pe_101
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[100]),
    .conf_bus_in(conf_bus_100),
    .branch_in(net_branch2peb_100),
    .branch_out(pe2net_branch_100),
    .ina(net2pea_100),
    .inb(net2peb_100),
    .outa(pe2neta_100),
    .outb(pe2netb_100)
  );


  cgra0_pe
  #(
    .PE_ID(102)
  )
  pe_102
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[101]),
    .conf_bus_in(conf_bus_101),
    .branch_in(net_branch2peb_101),
    .branch_out(pe2net_branch_101),
    .ina(net2pea_101),
    .inb(net2peb_101),
    .outa(pe2neta_101),
    .outb(pe2netb_101)
  );


  cgra0_pe
  #(
    .PE_ID(103)
  )
  pe_103
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[102]),
    .conf_bus_in(conf_bus_102),
    .branch_in(net_branch2peb_102),
    .branch_out(pe2net_branch_102),
    .ina(net2pea_102),
    .inb(net2peb_102),
    .outa(pe2neta_102),
    .outb(pe2netb_102)
  );


  cgra0_pe
  #(
    .PE_ID(104)
  )
  pe_104
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[103]),
    .conf_bus_in(conf_bus_103),
    .branch_in(net_branch2peb_103),
    .branch_out(pe2net_branch_103),
    .ina(net2pea_103),
    .inb(net2peb_103),
    .outa(pe2neta_103),
    .outb(pe2netb_103)
  );


  cgra0_pe
  #(
    .PE_ID(105)
  )
  pe_105
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[104]),
    .conf_bus_in(conf_bus_104),
    .branch_in(net_branch2peb_104),
    .branch_out(pe2net_branch_104),
    .ina(net2pea_104),
    .inb(net2peb_104),
    .outa(pe2neta_104),
    .outb(pe2netb_104)
  );


  cgra0_pe
  #(
    .PE_ID(106)
  )
  pe_106
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[105]),
    .conf_bus_in(conf_bus_105),
    .branch_in(net_branch2peb_105),
    .branch_out(pe2net_branch_105),
    .ina(net2pea_105),
    .inb(net2peb_105),
    .outa(pe2neta_105),
    .outb(pe2netb_105)
  );


  cgra0_pe
  #(
    .PE_ID(107)
  )
  pe_107
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[106]),
    .conf_bus_in(conf_bus_106),
    .branch_in(net_branch2peb_106),
    .branch_out(pe2net_branch_106),
    .ina(net2pea_106),
    .inb(net2peb_106),
    .outa(pe2neta_106),
    .outb(pe2netb_106)
  );


  cgra0_pe
  #(
    .PE_ID(108)
  )
  pe_108
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[107]),
    .conf_bus_in(conf_bus_107),
    .branch_in(net_branch2peb_107),
    .branch_out(pe2net_branch_107),
    .ina(net2pea_107),
    .inb(net2peb_107),
    .outa(pe2neta_107),
    .outb(pe2netb_107)
  );


  cgra0_pe
  #(
    .PE_ID(109)
  )
  pe_109
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[108]),
    .conf_bus_in(conf_bus_108),
    .branch_in(net_branch2peb_108),
    .branch_out(pe2net_branch_108),
    .ina(net2pea_108),
    .inb(net2peb_108),
    .outa(pe2neta_108),
    .outb(pe2netb_108)
  );


  cgra0_pe
  #(
    .PE_ID(110)
  )
  pe_110
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[109]),
    .conf_bus_in(conf_bus_109),
    .branch_in(net_branch2peb_109),
    .branch_out(pe2net_branch_109),
    .ina(net2pea_109),
    .inb(net2peb_109),
    .outa(pe2neta_109),
    .outb(pe2netb_109)
  );


  cgra0_pe
  #(
    .PE_ID(111)
  )
  pe_111
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[110]),
    .conf_bus_in(conf_bus_110),
    .branch_in(net_branch2peb_110),
    .branch_out(pe2net_branch_110),
    .ina(net2pea_110),
    .inb(net2peb_110),
    .outa(pe2neta_110),
    .outb(pe2netb_110)
  );


  cgra0_pe
  #(
    .PE_ID(112)
  )
  pe_112
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[111]),
    .conf_bus_in(conf_bus_111),
    .branch_in(net_branch2peb_111),
    .branch_out(pe2net_branch_111),
    .ina(net2pea_111),
    .inb(net2peb_111),
    .outa(pe2neta_111),
    .outb(pe2netb_111)
  );


  cgra0_pe
  #(
    .PE_ID(113)
  )
  pe_113
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[112]),
    .conf_bus_in(conf_bus_112),
    .branch_in(net_branch2peb_112),
    .branch_out(pe2net_branch_112),
    .ina(net2pea_112),
    .inb(net2peb_112),
    .outa(pe2neta_112),
    .outb(pe2netb_112)
  );


  cgra0_pe
  #(
    .PE_ID(114)
  )
  pe_114
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[113]),
    .conf_bus_in(conf_bus_113),
    .branch_in(net_branch2peb_113),
    .branch_out(pe2net_branch_113),
    .ina(net2pea_113),
    .inb(net2peb_113),
    .outa(pe2neta_113),
    .outb(pe2netb_113)
  );


  cgra0_pe
  #(
    .PE_ID(115)
  )
  pe_115
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[114]),
    .conf_bus_in(conf_bus_114),
    .branch_in(net_branch2peb_114),
    .branch_out(pe2net_branch_114),
    .ina(net2pea_114),
    .inb(net2peb_114),
    .outa(pe2neta_114),
    .outb(pe2netb_114)
  );


  cgra0_pe
  #(
    .PE_ID(116)
  )
  pe_116
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[115]),
    .conf_bus_in(conf_bus_115),
    .branch_in(net_branch2peb_115),
    .branch_out(pe2net_branch_115),
    .ina(net2pea_115),
    .inb(net2peb_115),
    .outa(pe2neta_115),
    .outb(pe2netb_115)
  );


  cgra0_pe
  #(
    .PE_ID(117)
  )
  pe_117
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[116]),
    .conf_bus_in(conf_bus_116),
    .branch_in(net_branch2peb_116),
    .branch_out(pe2net_branch_116),
    .ina(net2pea_116),
    .inb(net2peb_116),
    .outa(pe2neta_116),
    .outb(pe2netb_116)
  );


  cgra0_pe
  #(
    .PE_ID(118)
  )
  pe_118
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[117]),
    .conf_bus_in(conf_bus_117),
    .branch_in(net_branch2peb_117),
    .branch_out(pe2net_branch_117),
    .ina(net2pea_117),
    .inb(net2peb_117),
    .outa(pe2neta_117),
    .outb(pe2netb_117)
  );


  cgra0_pe
  #(
    .PE_ID(119)
  )
  pe_119
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[118]),
    .conf_bus_in(conf_bus_118),
    .branch_in(net_branch2peb_118),
    .branch_out(pe2net_branch_118),
    .ina(net2pea_118),
    .inb(net2peb_118),
    .outa(pe2neta_118),
    .outb(pe2netb_118)
  );


  cgra0_pe
  #(
    .PE_ID(120)
  )
  pe_120
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[119]),
    .conf_bus_in(conf_bus_119),
    .branch_in(net_branch2peb_119),
    .branch_out(pe2net_branch_119),
    .ina(net2pea_119),
    .inb(net2peb_119),
    .outa(pe2neta_119),
    .outb(pe2netb_119)
  );


  cgra0_pe
  #(
    .PE_ID(121)
  )
  pe_121
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[120]),
    .conf_bus_in(conf_bus_120),
    .branch_in(net_branch2peb_120),
    .branch_out(pe2net_branch_120),
    .ina(net2pea_120),
    .inb(net2peb_120),
    .outa(pe2neta_120),
    .outb(pe2netb_120)
  );


  cgra0_pe
  #(
    .PE_ID(122)
  )
  pe_122
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[121]),
    .conf_bus_in(conf_bus_121),
    .branch_in(net_branch2peb_121),
    .branch_out(pe2net_branch_121),
    .ina(net2pea_121),
    .inb(net2peb_121),
    .outa(pe2neta_121),
    .outb(pe2netb_121)
  );


  cgra0_pe
  #(
    .PE_ID(123)
  )
  pe_123
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[122]),
    .conf_bus_in(conf_bus_122),
    .branch_in(net_branch2peb_122),
    .branch_out(pe2net_branch_122),
    .ina(net2pea_122),
    .inb(net2peb_122),
    .outa(pe2neta_122),
    .outb(pe2netb_122)
  );


  cgra0_pe
  #(
    .PE_ID(124)
  )
  pe_124
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[123]),
    .conf_bus_in(conf_bus_123),
    .branch_in(net_branch2peb_123),
    .branch_out(pe2net_branch_123),
    .ina(net2pea_123),
    .inb(net2peb_123),
    .outa(pe2neta_123),
    .outb(pe2netb_123)
  );


  cgra0_pe
  #(
    .PE_ID(125)
  )
  pe_125
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[124]),
    .conf_bus_in(conf_bus_124),
    .branch_in(net_branch2peb_124),
    .branch_out(pe2net_branch_124),
    .ina(net2pea_124),
    .inb(net2peb_124),
    .outa(pe2neta_124),
    .outb(pe2netb_124)
  );


  cgra0_pe
  #(
    .PE_ID(126)
  )
  pe_126
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[125]),
    .conf_bus_in(conf_bus_125),
    .branch_in(net_branch2peb_125),
    .branch_out(pe2net_branch_125),
    .ina(net2pea_125),
    .inb(net2peb_125),
    .outa(pe2neta_125),
    .outb(pe2netb_125)
  );


  cgra0_pe
  #(
    .PE_ID(127)
  )
  pe_127
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[126]),
    .conf_bus_in(conf_bus_126),
    .branch_in(net_branch2peb_126),
    .branch_out(pe2net_branch_126),
    .ina(net2pea_126),
    .inb(net2peb_126),
    .outa(pe2neta_126),
    .outb(pe2netb_126)
  );


  cgra0_pe
  #(
    .PE_ID(128)
  )
  pe_128
  (
    .clk(clk),
    .rst(rst),
    .en(pes_en[127]),
    .conf_bus_in(conf_bus_127),
    .branch_in(net_branch2peb_127),
    .branch_out(pe2net_branch_127),
    .ina(net2pea_127),
    .inb(net2peb_127),
    .outa(pe2neta_127),
    .outb(pe2netb_127)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_0),
    .out(conf_bus_1)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_1),
    .out(conf_bus_2)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_2),
    .out(conf_bus_3)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_3),
    .out(conf_bus_4)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_4),
    .out(conf_bus_5)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_5),
    .out(conf_bus_6)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_6),
    .out(conf_bus_7)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_7),
    .out(conf_bus_8)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_8),
    .out(conf_bus_9)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_9),
    .out(conf_bus_10)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_10),
    .out(conf_bus_11)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_11),
    .out(conf_bus_12)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_12),
    .out(conf_bus_13)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_13),
    .out(conf_bus_14)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_14),
    .out(conf_bus_15)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_15),
    .out(conf_bus_16)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_16),
    .out(conf_bus_17)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_17),
    .out(conf_bus_18)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_18),
    .out(conf_bus_19)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_19),
    .out(conf_bus_20)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_20),
    .out(conf_bus_21)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_21),
    .out(conf_bus_22)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_22),
    .out(conf_bus_23)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_23),
    .out(conf_bus_24)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_24),
    .out(conf_bus_25)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_25),
    .out(conf_bus_26)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_26),
    .out(conf_bus_27)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_27),
    .out(conf_bus_28)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_28),
    .out(conf_bus_29)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_29),
    .out(conf_bus_30)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_30),
    .out(conf_bus_31)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_31),
    .out(conf_bus_32)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_32),
    .out(conf_bus_33)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_33),
    .out(conf_bus_34)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_34),
    .out(conf_bus_35)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_35),
    .out(conf_bus_36)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_36),
    .out(conf_bus_37)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_37),
    .out(conf_bus_38)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_38),
    .out(conf_bus_39)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_39),
    .out(conf_bus_40)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_40),
    .out(conf_bus_41)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_41),
    .out(conf_bus_42)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_42),
    .out(conf_bus_43)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_43),
    .out(conf_bus_44)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_44),
    .out(conf_bus_45)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_45),
    .out(conf_bus_46)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_46),
    .out(conf_bus_47)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_47),
    .out(conf_bus_48)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_48),
    .out(conf_bus_49)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_49),
    .out(conf_bus_50)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_50),
    .out(conf_bus_51)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_51),
    .out(conf_bus_52)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_52),
    .out(conf_bus_53)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_53),
    .out(conf_bus_54)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_54),
    .out(conf_bus_55)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_55),
    .out(conf_bus_56)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_56),
    .out(conf_bus_57)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_57),
    .out(conf_bus_58)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_58),
    .out(conf_bus_59)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_59),
    .out(conf_bus_60)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_60),
    .out(conf_bus_61)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_61),
    .out(conf_bus_62)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_62),
    .out(conf_bus_63)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_63),
    .out(conf_bus_64)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_64),
    .out(conf_bus_65)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_65),
    .out(conf_bus_66)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_66),
    .out(conf_bus_67)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_67),
    .out(conf_bus_68)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_68),
    .out(conf_bus_69)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_69),
    .out(conf_bus_70)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_70),
    .out(conf_bus_71)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_71),
    .out(conf_bus_72)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_72),
    .out(conf_bus_73)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_73),
    .out(conf_bus_74)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_74),
    .out(conf_bus_75)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_75),
    .out(conf_bus_76)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_76),
    .out(conf_bus_77)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_77),
    .out(conf_bus_78)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_78),
    .out(conf_bus_79)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_79),
    .out(conf_bus_80)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_80),
    .out(conf_bus_81)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_81),
    .out(conf_bus_82)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_82),
    .out(conf_bus_83)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_83),
    .out(conf_bus_84)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_84),
    .out(conf_bus_85)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_85),
    .out(conf_bus_86)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_86),
    .out(conf_bus_87)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_87),
    .out(conf_bus_88)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_88),
    .out(conf_bus_89)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_89),
    .out(conf_bus_90)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_90),
    .out(conf_bus_91)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_91),
    .out(conf_bus_92)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_92),
    .out(conf_bus_93)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_93),
    .out(conf_bus_94)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_94),
    .out(conf_bus_95)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_95),
    .out(conf_bus_96)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_96),
    .out(conf_bus_97)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_97),
    .out(conf_bus_98)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_98),
    .out(conf_bus_99)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_99),
    .out(conf_bus_100)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_100),
    .out(conf_bus_101)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_101),
    .out(conf_bus_102)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_102),
    .out(conf_bus_103)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_103),
    .out(conf_bus_104)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_104),
    .out(conf_bus_105)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_105),
    .out(conf_bus_106)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_106),
    .out(conf_bus_107)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_107),
    .out(conf_bus_108)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_108),
    .out(conf_bus_109)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_109),
    .out(conf_bus_110)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_110),
    .out(conf_bus_111)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_111),
    .out(conf_bus_112)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_112),
    .out(conf_bus_113)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_113),
    .out(conf_bus_114)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_114),
    .out(conf_bus_115)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_115),
    .out(conf_bus_116)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_116),
    .out(conf_bus_117)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_117),
    .out(conf_bus_118)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_118),
    .out(conf_bus_119)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_119),
    .out(conf_bus_120)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_120),
    .out(conf_bus_121)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_121),
    .out(conf_bus_122)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_122),
    .out(conf_bus_123)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_123),
    .out(conf_bus_124)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_124),
    .out(conf_bus_125)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_125),
    .out(conf_bus_126)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_126),
    .out(conf_bus_127)
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_127),
    .out(conf_bus_128)
  );


  omega256x256_4_0_8
  #(
    .WIDTH(16),
    .PIPE_EXTRA(0)
  )
  net
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net),
    .en(net_en),
    .net_conf_bus_in(conf_bus_128),
    .in0(pe2neta_0),
    .in1(pe2netb_0),
    .in2(pe2neta_1),
    .in3(pe2netb_1),
    .in4(pe2neta_2),
    .in5(pe2netb_2),
    .in6(pe2neta_3),
    .in7(pe2netb_3),
    .in8(pe2neta_4),
    .in9(pe2netb_4),
    .in10(pe2neta_5),
    .in11(pe2netb_5),
    .in12(pe2neta_6),
    .in13(pe2netb_6),
    .in14(pe2neta_7),
    .in15(pe2netb_7),
    .in16(pe2neta_8),
    .in17(pe2netb_8),
    .in18(pe2neta_9),
    .in19(pe2netb_9),
    .in20(pe2neta_10),
    .in21(pe2netb_10),
    .in22(pe2neta_11),
    .in23(pe2netb_11),
    .in24(pe2neta_12),
    .in25(pe2netb_12),
    .in26(pe2neta_13),
    .in27(pe2netb_13),
    .in28(pe2neta_14),
    .in29(pe2netb_14),
    .in30(pe2neta_15),
    .in31(pe2netb_15),
    .in32(pe2neta_16),
    .in33(pe2netb_16),
    .in34(pe2neta_17),
    .in35(pe2netb_17),
    .in36(pe2neta_18),
    .in37(pe2netb_18),
    .in38(pe2neta_19),
    .in39(pe2netb_19),
    .in40(pe2neta_20),
    .in41(pe2netb_20),
    .in42(pe2neta_21),
    .in43(pe2netb_21),
    .in44(pe2neta_22),
    .in45(pe2netb_22),
    .in46(pe2neta_23),
    .in47(pe2netb_23),
    .in48(pe2neta_24),
    .in49(pe2netb_24),
    .in50(pe2neta_25),
    .in51(pe2netb_25),
    .in52(pe2neta_26),
    .in53(pe2netb_26),
    .in54(pe2neta_27),
    .in55(pe2netb_27),
    .in56(pe2neta_28),
    .in57(pe2netb_28),
    .in58(pe2neta_29),
    .in59(pe2netb_29),
    .in60(pe2neta_30),
    .in61(pe2netb_30),
    .in62(pe2neta_31),
    .in63(pe2netb_31),
    .in64(pe2neta_32),
    .in65(pe2netb_32),
    .in66(pe2neta_33),
    .in67(pe2netb_33),
    .in68(pe2neta_34),
    .in69(pe2netb_34),
    .in70(pe2neta_35),
    .in71(pe2netb_35),
    .in72(pe2neta_36),
    .in73(pe2netb_36),
    .in74(pe2neta_37),
    .in75(pe2netb_37),
    .in76(pe2neta_38),
    .in77(pe2netb_38),
    .in78(pe2neta_39),
    .in79(pe2netb_39),
    .in80(pe2neta_40),
    .in81(pe2netb_40),
    .in82(pe2neta_41),
    .in83(pe2netb_41),
    .in84(pe2neta_42),
    .in85(pe2netb_42),
    .in86(pe2neta_43),
    .in87(pe2netb_43),
    .in88(pe2neta_44),
    .in89(pe2netb_44),
    .in90(pe2neta_45),
    .in91(pe2netb_45),
    .in92(pe2neta_46),
    .in93(pe2netb_46),
    .in94(pe2neta_47),
    .in95(pe2netb_47),
    .in96(pe2neta_48),
    .in97(pe2netb_48),
    .in98(pe2neta_49),
    .in99(pe2netb_49),
    .in100(pe2neta_50),
    .in101(pe2netb_50),
    .in102(pe2neta_51),
    .in103(pe2netb_51),
    .in104(pe2neta_52),
    .in105(pe2netb_52),
    .in106(pe2neta_53),
    .in107(pe2netb_53),
    .in108(pe2neta_54),
    .in109(pe2netb_54),
    .in110(pe2neta_55),
    .in111(pe2netb_55),
    .in112(pe2neta_56),
    .in113(pe2netb_56),
    .in114(pe2neta_57),
    .in115(pe2netb_57),
    .in116(pe2neta_58),
    .in117(pe2netb_58),
    .in118(pe2neta_59),
    .in119(pe2netb_59),
    .in120(pe2neta_60),
    .in121(pe2netb_60),
    .in122(pe2neta_61),
    .in123(pe2netb_61),
    .in124(pe2neta_62),
    .in125(pe2netb_62),
    .in126(pe2neta_63),
    .in127(pe2netb_63),
    .in128(pe2neta_64),
    .in129(pe2netb_64),
    .in130(pe2neta_65),
    .in131(pe2netb_65),
    .in132(pe2neta_66),
    .in133(pe2netb_66),
    .in134(pe2neta_67),
    .in135(pe2netb_67),
    .in136(pe2neta_68),
    .in137(pe2netb_68),
    .in138(pe2neta_69),
    .in139(pe2netb_69),
    .in140(pe2neta_70),
    .in141(pe2netb_70),
    .in142(pe2neta_71),
    .in143(pe2netb_71),
    .in144(pe2neta_72),
    .in145(pe2netb_72),
    .in146(pe2neta_73),
    .in147(pe2netb_73),
    .in148(pe2neta_74),
    .in149(pe2netb_74),
    .in150(pe2neta_75),
    .in151(pe2netb_75),
    .in152(pe2neta_76),
    .in153(pe2netb_76),
    .in154(pe2neta_77),
    .in155(pe2netb_77),
    .in156(pe2neta_78),
    .in157(pe2netb_78),
    .in158(pe2neta_79),
    .in159(pe2netb_79),
    .in160(pe2neta_80),
    .in161(pe2netb_80),
    .in162(pe2neta_81),
    .in163(pe2netb_81),
    .in164(pe2neta_82),
    .in165(pe2netb_82),
    .in166(pe2neta_83),
    .in167(pe2netb_83),
    .in168(pe2neta_84),
    .in169(pe2netb_84),
    .in170(pe2neta_85),
    .in171(pe2netb_85),
    .in172(pe2neta_86),
    .in173(pe2netb_86),
    .in174(pe2neta_87),
    .in175(pe2netb_87),
    .in176(pe2neta_88),
    .in177(pe2netb_88),
    .in178(pe2neta_89),
    .in179(pe2netb_89),
    .in180(pe2neta_90),
    .in181(pe2netb_90),
    .in182(pe2neta_91),
    .in183(pe2netb_91),
    .in184(pe2neta_92),
    .in185(pe2netb_92),
    .in186(pe2neta_93),
    .in187(pe2netb_93),
    .in188(pe2neta_94),
    .in189(pe2netb_94),
    .in190(pe2neta_95),
    .in191(pe2netb_95),
    .in192(pe2neta_96),
    .in193(pe2netb_96),
    .in194(pe2neta_97),
    .in195(pe2netb_97),
    .in196(pe2neta_98),
    .in197(pe2netb_98),
    .in198(pe2neta_99),
    .in199(pe2netb_99),
    .in200(pe2neta_100),
    .in201(pe2netb_100),
    .in202(pe2neta_101),
    .in203(pe2netb_101),
    .in204(pe2neta_102),
    .in205(pe2netb_102),
    .in206(pe2neta_103),
    .in207(pe2netb_103),
    .in208(pe2neta_104),
    .in209(pe2netb_104),
    .in210(pe2neta_105),
    .in211(pe2netb_105),
    .in212(pe2neta_106),
    .in213(pe2netb_106),
    .in214(pe2neta_107),
    .in215(pe2netb_107),
    .in216(pe2neta_108),
    .in217(pe2netb_108),
    .in218(pe2neta_109),
    .in219(pe2netb_109),
    .in220(pe2neta_110),
    .in221(pe2netb_110),
    .in222(pe2neta_111),
    .in223(pe2netb_111),
    .in224(pe2neta_112),
    .in225(pe2netb_112),
    .in226(pe2neta_113),
    .in227(pe2netb_113),
    .in228(pe2neta_114),
    .in229(pe2netb_114),
    .in230(pe2neta_115),
    .in231(pe2netb_115),
    .in232(pe2neta_116),
    .in233(pe2netb_116),
    .in234(pe2neta_117),
    .in235(pe2netb_117),
    .in236(pe2neta_118),
    .in237(pe2netb_118),
    .in238(pe2neta_119),
    .in239(pe2netb_119),
    .in240(pe2neta_120),
    .in241(pe2netb_120),
    .in242(pe2neta_121),
    .in243(pe2netb_121),
    .in244(pe2neta_122),
    .in245(pe2netb_122),
    .in246(pe2neta_123),
    .in247(pe2netb_123),
    .in248(pe2neta_124),
    .in249(pe2netb_124),
    .in250(pe2neta_125),
    .in251(pe2netb_125),
    .in252(pe2neta_126),
    .in253(pe2netb_126),
    .in254(pe2neta_127),
    .in255(pe2netb_127),
    .out0(net2pea_0),
    .out1(net2peb_0),
    .out2(net2pea_1),
    .out3(net2peb_1),
    .out4(net2pea_2),
    .out5(net2peb_2),
    .out6(net2pea_3),
    .out7(net2peb_3),
    .out8(net2pea_4),
    .out9(net2peb_4),
    .out10(net2pea_5),
    .out11(net2peb_5),
    .out12(net2pea_6),
    .out13(net2peb_6),
    .out14(net2pea_7),
    .out15(net2peb_7),
    .out16(net2pea_8),
    .out17(net2peb_8),
    .out18(net2pea_9),
    .out19(net2peb_9),
    .out20(net2pea_10),
    .out21(net2peb_10),
    .out22(net2pea_11),
    .out23(net2peb_11),
    .out24(net2pea_12),
    .out25(net2peb_12),
    .out26(net2pea_13),
    .out27(net2peb_13),
    .out28(net2pea_14),
    .out29(net2peb_14),
    .out30(net2pea_15),
    .out31(net2peb_15),
    .out32(net2pea_16),
    .out33(net2peb_16),
    .out34(net2pea_17),
    .out35(net2peb_17),
    .out36(net2pea_18),
    .out37(net2peb_18),
    .out38(net2pea_19),
    .out39(net2peb_19),
    .out40(net2pea_20),
    .out41(net2peb_20),
    .out42(net2pea_21),
    .out43(net2peb_21),
    .out44(net2pea_22),
    .out45(net2peb_22),
    .out46(net2pea_23),
    .out47(net2peb_23),
    .out48(net2pea_24),
    .out49(net2peb_24),
    .out50(net2pea_25),
    .out51(net2peb_25),
    .out52(net2pea_26),
    .out53(net2peb_26),
    .out54(net2pea_27),
    .out55(net2peb_27),
    .out56(net2pea_28),
    .out57(net2peb_28),
    .out58(net2pea_29),
    .out59(net2peb_29),
    .out60(net2pea_30),
    .out61(net2peb_30),
    .out62(net2pea_31),
    .out63(net2peb_31),
    .out64(net2pea_32),
    .out65(net2peb_32),
    .out66(net2pea_33),
    .out67(net2peb_33),
    .out68(net2pea_34),
    .out69(net2peb_34),
    .out70(net2pea_35),
    .out71(net2peb_35),
    .out72(net2pea_36),
    .out73(net2peb_36),
    .out74(net2pea_37),
    .out75(net2peb_37),
    .out76(net2pea_38),
    .out77(net2peb_38),
    .out78(net2pea_39),
    .out79(net2peb_39),
    .out80(net2pea_40),
    .out81(net2peb_40),
    .out82(net2pea_41),
    .out83(net2peb_41),
    .out84(net2pea_42),
    .out85(net2peb_42),
    .out86(net2pea_43),
    .out87(net2peb_43),
    .out88(net2pea_44),
    .out89(net2peb_44),
    .out90(net2pea_45),
    .out91(net2peb_45),
    .out92(net2pea_46),
    .out93(net2peb_46),
    .out94(net2pea_47),
    .out95(net2peb_47),
    .out96(net2pea_48),
    .out97(net2peb_48),
    .out98(net2pea_49),
    .out99(net2peb_49),
    .out100(net2pea_50),
    .out101(net2peb_50),
    .out102(net2pea_51),
    .out103(net2peb_51),
    .out104(net2pea_52),
    .out105(net2peb_52),
    .out106(net2pea_53),
    .out107(net2peb_53),
    .out108(net2pea_54),
    .out109(net2peb_54),
    .out110(net2pea_55),
    .out111(net2peb_55),
    .out112(net2pea_56),
    .out113(net2peb_56),
    .out114(net2pea_57),
    .out115(net2peb_57),
    .out116(net2pea_58),
    .out117(net2peb_58),
    .out118(net2pea_59),
    .out119(net2peb_59),
    .out120(net2pea_60),
    .out121(net2peb_60),
    .out122(net2pea_61),
    .out123(net2peb_61),
    .out124(net2pea_62),
    .out125(net2peb_62),
    .out126(net2pea_63),
    .out127(net2peb_63),
    .out128(net2pea_64),
    .out129(net2peb_64),
    .out130(net2pea_65),
    .out131(net2peb_65),
    .out132(net2pea_66),
    .out133(net2peb_66),
    .out134(net2pea_67),
    .out135(net2peb_67),
    .out136(net2pea_68),
    .out137(net2peb_68),
    .out138(net2pea_69),
    .out139(net2peb_69),
    .out140(net2pea_70),
    .out141(net2peb_70),
    .out142(net2pea_71),
    .out143(net2peb_71),
    .out144(net2pea_72),
    .out145(net2peb_72),
    .out146(net2pea_73),
    .out147(net2peb_73),
    .out148(net2pea_74),
    .out149(net2peb_74),
    .out150(net2pea_75),
    .out151(net2peb_75),
    .out152(net2pea_76),
    .out153(net2peb_76),
    .out154(net2pea_77),
    .out155(net2peb_77),
    .out156(net2pea_78),
    .out157(net2peb_78),
    .out158(net2pea_79),
    .out159(net2peb_79),
    .out160(net2pea_80),
    .out161(net2peb_80),
    .out162(net2pea_81),
    .out163(net2peb_81),
    .out164(net2pea_82),
    .out165(net2peb_82),
    .out166(net2pea_83),
    .out167(net2peb_83),
    .out168(net2pea_84),
    .out169(net2peb_84),
    .out170(net2pea_85),
    .out171(net2peb_85),
    .out172(net2pea_86),
    .out173(net2peb_86),
    .out174(net2pea_87),
    .out175(net2peb_87),
    .out176(net2pea_88),
    .out177(net2peb_88),
    .out178(net2pea_89),
    .out179(net2peb_89),
    .out180(net2pea_90),
    .out181(net2peb_90),
    .out182(net2pea_91),
    .out183(net2peb_91),
    .out184(net2pea_92),
    .out185(net2peb_92),
    .out186(net2pea_93),
    .out187(net2peb_93),
    .out188(net2pea_94),
    .out189(net2peb_94),
    .out190(net2pea_95),
    .out191(net2peb_95),
    .out192(net2pea_96),
    .out193(net2peb_96),
    .out194(net2pea_97),
    .out195(net2peb_97),
    .out196(net2pea_98),
    .out197(net2peb_98),
    .out198(net2pea_99),
    .out199(net2peb_99),
    .out200(net2pea_100),
    .out201(net2peb_100),
    .out202(net2pea_101),
    .out203(net2peb_101),
    .out204(net2pea_102),
    .out205(net2peb_102),
    .out206(net2pea_103),
    .out207(net2peb_103),
    .out208(net2pea_104),
    .out209(net2peb_104),
    .out210(net2pea_105),
    .out211(net2peb_105),
    .out212(net2pea_106),
    .out213(net2peb_106),
    .out214(net2pea_107),
    .out215(net2peb_107),
    .out216(net2pea_108),
    .out217(net2peb_108),
    .out218(net2pea_109),
    .out219(net2peb_109),
    .out220(net2pea_110),
    .out221(net2peb_110),
    .out222(net2pea_111),
    .out223(net2peb_111),
    .out224(net2pea_112),
    .out225(net2peb_112),
    .out226(net2pea_113),
    .out227(net2peb_113),
    .out228(net2pea_114),
    .out229(net2peb_114),
    .out230(net2pea_115),
    .out231(net2peb_115),
    .out232(net2pea_116),
    .out233(net2peb_116),
    .out234(net2pea_117),
    .out235(net2peb_117),
    .out236(net2pea_118),
    .out237(net2peb_118),
    .out238(net2pea_119),
    .out239(net2peb_119),
    .out240(net2pea_120),
    .out241(net2peb_120),
    .out242(net2pea_121),
    .out243(net2peb_121),
    .out244(net2pea_122),
    .out245(net2peb_122),
    .out246(net2pea_123),
    .out247(net2peb_123),
    .out248(net2pea_124),
    .out249(net2peb_124),
    .out250(net2pea_125),
    .out251(net2peb_125),
    .out252(net2pea_126),
    .out253(net2peb_126),
    .out254(net2pea_127),
    .out255(net2peb_127)
  );


  omega_branch128x128_4_0_8
  #(
    .WIDTH(1),
    .PIPE_EXTRA(0)
  )
  net_branch
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[127:0]),
    .en(net_en[639:0]),
    .net_conf_bus_in(conf_bus_128),
    .in0(pe2net_branch_0),
    .in1(pe2net_branch_1),
    .in2(pe2net_branch_2),
    .in3(pe2net_branch_3),
    .in4(pe2net_branch_4),
    .in5(pe2net_branch_5),
    .in6(pe2net_branch_6),
    .in7(pe2net_branch_7),
    .in8(pe2net_branch_8),
    .in9(pe2net_branch_9),
    .in10(pe2net_branch_10),
    .in11(pe2net_branch_11),
    .in12(pe2net_branch_12),
    .in13(pe2net_branch_13),
    .in14(pe2net_branch_14),
    .in15(pe2net_branch_15),
    .in16(pe2net_branch_16),
    .in17(pe2net_branch_17),
    .in18(pe2net_branch_18),
    .in19(pe2net_branch_19),
    .in20(pe2net_branch_20),
    .in21(pe2net_branch_21),
    .in22(pe2net_branch_22),
    .in23(pe2net_branch_23),
    .in24(pe2net_branch_24),
    .in25(pe2net_branch_25),
    .in26(pe2net_branch_26),
    .in27(pe2net_branch_27),
    .in28(pe2net_branch_28),
    .in29(pe2net_branch_29),
    .in30(pe2net_branch_30),
    .in31(pe2net_branch_31),
    .in32(pe2net_branch_32),
    .in33(pe2net_branch_33),
    .in34(pe2net_branch_34),
    .in35(pe2net_branch_35),
    .in36(pe2net_branch_36),
    .in37(pe2net_branch_37),
    .in38(pe2net_branch_38),
    .in39(pe2net_branch_39),
    .in40(pe2net_branch_40),
    .in41(pe2net_branch_41),
    .in42(pe2net_branch_42),
    .in43(pe2net_branch_43),
    .in44(pe2net_branch_44),
    .in45(pe2net_branch_45),
    .in46(pe2net_branch_46),
    .in47(pe2net_branch_47),
    .in48(pe2net_branch_48),
    .in49(pe2net_branch_49),
    .in50(pe2net_branch_50),
    .in51(pe2net_branch_51),
    .in52(pe2net_branch_52),
    .in53(pe2net_branch_53),
    .in54(pe2net_branch_54),
    .in55(pe2net_branch_55),
    .in56(pe2net_branch_56),
    .in57(pe2net_branch_57),
    .in58(pe2net_branch_58),
    .in59(pe2net_branch_59),
    .in60(pe2net_branch_60),
    .in61(pe2net_branch_61),
    .in62(pe2net_branch_62),
    .in63(pe2net_branch_63),
    .in64(pe2net_branch_64),
    .in65(pe2net_branch_65),
    .in66(pe2net_branch_66),
    .in67(pe2net_branch_67),
    .in68(pe2net_branch_68),
    .in69(pe2net_branch_69),
    .in70(pe2net_branch_70),
    .in71(pe2net_branch_71),
    .in72(pe2net_branch_72),
    .in73(pe2net_branch_73),
    .in74(pe2net_branch_74),
    .in75(pe2net_branch_75),
    .in76(pe2net_branch_76),
    .in77(pe2net_branch_77),
    .in78(pe2net_branch_78),
    .in79(pe2net_branch_79),
    .in80(pe2net_branch_80),
    .in81(pe2net_branch_81),
    .in82(pe2net_branch_82),
    .in83(pe2net_branch_83),
    .in84(pe2net_branch_84),
    .in85(pe2net_branch_85),
    .in86(pe2net_branch_86),
    .in87(pe2net_branch_87),
    .in88(pe2net_branch_88),
    .in89(pe2net_branch_89),
    .in90(pe2net_branch_90),
    .in91(pe2net_branch_91),
    .in92(pe2net_branch_92),
    .in93(pe2net_branch_93),
    .in94(pe2net_branch_94),
    .in95(pe2net_branch_95),
    .in96(pe2net_branch_96),
    .in97(pe2net_branch_97),
    .in98(pe2net_branch_98),
    .in99(pe2net_branch_99),
    .in100(pe2net_branch_100),
    .in101(pe2net_branch_101),
    .in102(pe2net_branch_102),
    .in103(pe2net_branch_103),
    .in104(pe2net_branch_104),
    .in105(pe2net_branch_105),
    .in106(pe2net_branch_106),
    .in107(pe2net_branch_107),
    .in108(pe2net_branch_108),
    .in109(pe2net_branch_109),
    .in110(pe2net_branch_110),
    .in111(pe2net_branch_111),
    .in112(pe2net_branch_112),
    .in113(pe2net_branch_113),
    .in114(pe2net_branch_114),
    .in115(pe2net_branch_115),
    .in116(pe2net_branch_116),
    .in117(pe2net_branch_117),
    .in118(pe2net_branch_118),
    .in119(pe2net_branch_119),
    .in120(pe2net_branch_120),
    .in121(pe2net_branch_121),
    .in122(pe2net_branch_122),
    .in123(pe2net_branch_123),
    .in124(pe2net_branch_124),
    .in125(pe2net_branch_125),
    .in126(pe2net_branch_126),
    .in127(pe2net_branch_127),
    .out0(net_branch2peb_0),
    .out1(net_branch2peb_1),
    .out2(net_branch2peb_2),
    .out3(net_branch2peb_3),
    .out4(net_branch2peb_4),
    .out5(net_branch2peb_5),
    .out6(net_branch2peb_6),
    .out7(net_branch2peb_7),
    .out8(net_branch2peb_8),
    .out9(net_branch2peb_9),
    .out10(net_branch2peb_10),
    .out11(net_branch2peb_11),
    .out12(net_branch2peb_12),
    .out13(net_branch2peb_13),
    .out14(net_branch2peb_14),
    .out15(net_branch2peb_15),
    .out16(net_branch2peb_16),
    .out17(net_branch2peb_17),
    .out18(net_branch2peb_18),
    .out19(net_branch2peb_19),
    .out20(net_branch2peb_20),
    .out21(net_branch2peb_21),
    .out22(net_branch2peb_22),
    .out23(net_branch2peb_23),
    .out24(net_branch2peb_24),
    .out25(net_branch2peb_25),
    .out26(net_branch2peb_26),
    .out27(net_branch2peb_27),
    .out28(net_branch2peb_28),
    .out29(net_branch2peb_29),
    .out30(net_branch2peb_30),
    .out31(net_branch2peb_31),
    .out32(net_branch2peb_32),
    .out33(net_branch2peb_33),
    .out34(net_branch2peb_34),
    .out35(net_branch2peb_35),
    .out36(net_branch2peb_36),
    .out37(net_branch2peb_37),
    .out38(net_branch2peb_38),
    .out39(net_branch2peb_39),
    .out40(net_branch2peb_40),
    .out41(net_branch2peb_41),
    .out42(net_branch2peb_42),
    .out43(net_branch2peb_43),
    .out44(net_branch2peb_44),
    .out45(net_branch2peb_45),
    .out46(net_branch2peb_46),
    .out47(net_branch2peb_47),
    .out48(net_branch2peb_48),
    .out49(net_branch2peb_49),
    .out50(net_branch2peb_50),
    .out51(net_branch2peb_51),
    .out52(net_branch2peb_52),
    .out53(net_branch2peb_53),
    .out54(net_branch2peb_54),
    .out55(net_branch2peb_55),
    .out56(net_branch2peb_56),
    .out57(net_branch2peb_57),
    .out58(net_branch2peb_58),
    .out59(net_branch2peb_59),
    .out60(net_branch2peb_60),
    .out61(net_branch2peb_61),
    .out62(net_branch2peb_62),
    .out63(net_branch2peb_63),
    .out64(net_branch2peb_64),
    .out65(net_branch2peb_65),
    .out66(net_branch2peb_66),
    .out67(net_branch2peb_67),
    .out68(net_branch2peb_68),
    .out69(net_branch2peb_69),
    .out70(net_branch2peb_70),
    .out71(net_branch2peb_71),
    .out72(net_branch2peb_72),
    .out73(net_branch2peb_73),
    .out74(net_branch2peb_74),
    .out75(net_branch2peb_75),
    .out76(net_branch2peb_76),
    .out77(net_branch2peb_77),
    .out78(net_branch2peb_78),
    .out79(net_branch2peb_79),
    .out80(net_branch2peb_80),
    .out81(net_branch2peb_81),
    .out82(net_branch2peb_82),
    .out83(net_branch2peb_83),
    .out84(net_branch2peb_84),
    .out85(net_branch2peb_85),
    .out86(net_branch2peb_86),
    .out87(net_branch2peb_87),
    .out88(net_branch2peb_88),
    .out89(net_branch2peb_89),
    .out90(net_branch2peb_90),
    .out91(net_branch2peb_91),
    .out92(net_branch2peb_92),
    .out93(net_branch2peb_93),
    .out94(net_branch2peb_94),
    .out95(net_branch2peb_95),
    .out96(net_branch2peb_96),
    .out97(net_branch2peb_97),
    .out98(net_branch2peb_98),
    .out99(net_branch2peb_99),
    .out100(net_branch2peb_100),
    .out101(net_branch2peb_101),
    .out102(net_branch2peb_102),
    .out103(net_branch2peb_103),
    .out104(net_branch2peb_104),
    .out105(net_branch2peb_105),
    .out106(net_branch2peb_106),
    .out107(net_branch2peb_107),
    .out108(net_branch2peb_108),
    .out109(net_branch2peb_109),
    .out110(net_branch2peb_110),
    .out111(net_branch2peb_111),
    .out112(net_branch2peb_112),
    .out113(net_branch2peb_113),
    .out114(net_branch2peb_114),
    .out115(net_branch2peb_115),
    .out116(net_branch2peb_116),
    .out117(net_branch2peb_117),
    .out118(net_branch2peb_118),
    .out119(net_branch2peb_119),
    .out120(net_branch2peb_120),
    .out121(net_branch2peb_121),
    .out122(net_branch2peb_122),
    .out123(net_branch2peb_123),
    .out124(net_branch2peb_124),
    .out125(net_branch2peb_125),
    .out126(net_branch2peb_126),
    .out127(net_branch2peb_127)
  );

endmodule