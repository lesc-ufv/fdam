module cgra0_top
(
  input clk,
  input rst,
  input [128-1:0] pes_en,
  input [64-1:0] conf_bus_in,
  input [1280-1:0] net_en,
  input [256-1:0] en_pc_net,
  output [16-1:0] fifo_in_re,
  input [256-1:0] fifo_in_data,
  output [16-1:0] fifo_out_we,
  output [256-1:0] fifo_out_data
);


  wire [64-1:0] conf_bus [0:129-1];

  wire [16-1:0] pe2neta [0:128-1];
  wire [16-1:0] pe2netb [0:128-1];
  wire [16-1:0] net2pea [0:128-1];
  wire [16-1:0] net2peb [0:128-1];

  genvar genv;


  reg_pipe_
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  reg_conf_bus_in2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_in),
    .out(conf_bus[0])
  );


  generate for(genv=0; genv<16; genv=genv+1) begin : inst_pe_io

    cgra0_pe_io
    #(
      .PE_ID(genv + 1)
    )
    pe_io
    (
      .clk(clk),
      .rst(rst),
      .en(pes_en[genv]),
      .conf_bus_in(conf_bus[genv]),
      .fifo_in_re(fifo_in_re[genv]),
      .fifo_in_data(fifo_in_data[(genv+1)*16-1:genv*16]),
      .fifo_out_we(fifo_out_we[genv]),
      .fifo_out_data(fifo_out_data[(genv+1)*16-1:genv*16]),
      .ina(net2pea[genv]),
      .inb(net2peb[genv]),
      .outa(pe2neta[genv]),
      .outb(pe2netb[genv])
    );


    reg_pipe_
    #(
      .NUM_STAGES(1),
      .DATA_WIDTH(64)
    )
    conf_bus_reg_pe_io
    (
      .clk(clk),
      .rst(1'b0),
      .en(1'b1),
      .in(conf_bus[genv]),
      .out(conf_bus[genv + 1])
    );

  end
  endgenerate


  generate for(genv=16; genv<128; genv=genv+1) begin : inst_pe

    cgra0_pe
    #(
      .PE_ID(genv + 1)
    )
    pe
    (
      .clk(clk),
      .rst(rst),
      .en(pes_en[genv]),
      .conf_bus_in(conf_bus[genv]),
      .ina(net2pea[genv]),
      .inb(net2peb[genv]),
      .outa(pe2neta[genv]),
      .outb(pe2netb[genv])
    );


    reg_pipe_
    #(
      .NUM_STAGES(1),
      .DATA_WIDTH(64)
    )
    conf_bus_reg_pe
    (
      .clk(clk),
      .rst(1'b0),
      .en(1'b1),
      .in(conf_bus[genv]),
      .out(conf_bus[genv + 1])
    );

  end
  endgenerate


  omega256x256_4_0_8
  #(
    .WIDTH(16),
    .PIPE_EXTRA(0)
  )
  net
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net),
    .en(net_en),
    .net_conf_bus_in(conf_bus[128]),
    .in0(pe2neta[0]),
    .in1(pe2netb[0]),
    .in2(pe2neta[1]),
    .in3(pe2netb[1]),
    .in4(pe2neta[2]),
    .in5(pe2netb[2]),
    .in6(pe2neta[3]),
    .in7(pe2netb[3]),
    .in8(pe2neta[4]),
    .in9(pe2netb[4]),
    .in10(pe2neta[5]),
    .in11(pe2netb[5]),
    .in12(pe2neta[6]),
    .in13(pe2netb[6]),
    .in14(pe2neta[7]),
    .in15(pe2netb[7]),
    .in16(pe2neta[8]),
    .in17(pe2netb[8]),
    .in18(pe2neta[9]),
    .in19(pe2netb[9]),
    .in20(pe2neta[10]),
    .in21(pe2netb[10]),
    .in22(pe2neta[11]),
    .in23(pe2netb[11]),
    .in24(pe2neta[12]),
    .in25(pe2netb[12]),
    .in26(pe2neta[13]),
    .in27(pe2netb[13]),
    .in28(pe2neta[14]),
    .in29(pe2netb[14]),
    .in30(pe2neta[15]),
    .in31(pe2netb[15]),
    .in32(pe2neta[16]),
    .in33(pe2netb[16]),
    .in34(pe2neta[17]),
    .in35(pe2netb[17]),
    .in36(pe2neta[18]),
    .in37(pe2netb[18]),
    .in38(pe2neta[19]),
    .in39(pe2netb[19]),
    .in40(pe2neta[20]),
    .in41(pe2netb[20]),
    .in42(pe2neta[21]),
    .in43(pe2netb[21]),
    .in44(pe2neta[22]),
    .in45(pe2netb[22]),
    .in46(pe2neta[23]),
    .in47(pe2netb[23]),
    .in48(pe2neta[24]),
    .in49(pe2netb[24]),
    .in50(pe2neta[25]),
    .in51(pe2netb[25]),
    .in52(pe2neta[26]),
    .in53(pe2netb[26]),
    .in54(pe2neta[27]),
    .in55(pe2netb[27]),
    .in56(pe2neta[28]),
    .in57(pe2netb[28]),
    .in58(pe2neta[29]),
    .in59(pe2netb[29]),
    .in60(pe2neta[30]),
    .in61(pe2netb[30]),
    .in62(pe2neta[31]),
    .in63(pe2netb[31]),
    .in64(pe2neta[32]),
    .in65(pe2netb[32]),
    .in66(pe2neta[33]),
    .in67(pe2netb[33]),
    .in68(pe2neta[34]),
    .in69(pe2netb[34]),
    .in70(pe2neta[35]),
    .in71(pe2netb[35]),
    .in72(pe2neta[36]),
    .in73(pe2netb[36]),
    .in74(pe2neta[37]),
    .in75(pe2netb[37]),
    .in76(pe2neta[38]),
    .in77(pe2netb[38]),
    .in78(pe2neta[39]),
    .in79(pe2netb[39]),
    .in80(pe2neta[40]),
    .in81(pe2netb[40]),
    .in82(pe2neta[41]),
    .in83(pe2netb[41]),
    .in84(pe2neta[42]),
    .in85(pe2netb[42]),
    .in86(pe2neta[43]),
    .in87(pe2netb[43]),
    .in88(pe2neta[44]),
    .in89(pe2netb[44]),
    .in90(pe2neta[45]),
    .in91(pe2netb[45]),
    .in92(pe2neta[46]),
    .in93(pe2netb[46]),
    .in94(pe2neta[47]),
    .in95(pe2netb[47]),
    .in96(pe2neta[48]),
    .in97(pe2netb[48]),
    .in98(pe2neta[49]),
    .in99(pe2netb[49]),
    .in100(pe2neta[50]),
    .in101(pe2netb[50]),
    .in102(pe2neta[51]),
    .in103(pe2netb[51]),
    .in104(pe2neta[52]),
    .in105(pe2netb[52]),
    .in106(pe2neta[53]),
    .in107(pe2netb[53]),
    .in108(pe2neta[54]),
    .in109(pe2netb[54]),
    .in110(pe2neta[55]),
    .in111(pe2netb[55]),
    .in112(pe2neta[56]),
    .in113(pe2netb[56]),
    .in114(pe2neta[57]),
    .in115(pe2netb[57]),
    .in116(pe2neta[58]),
    .in117(pe2netb[58]),
    .in118(pe2neta[59]),
    .in119(pe2netb[59]),
    .in120(pe2neta[60]),
    .in121(pe2netb[60]),
    .in122(pe2neta[61]),
    .in123(pe2netb[61]),
    .in124(pe2neta[62]),
    .in125(pe2netb[62]),
    .in126(pe2neta[63]),
    .in127(pe2netb[63]),
    .in128(pe2neta[64]),
    .in129(pe2netb[64]),
    .in130(pe2neta[65]),
    .in131(pe2netb[65]),
    .in132(pe2neta[66]),
    .in133(pe2netb[66]),
    .in134(pe2neta[67]),
    .in135(pe2netb[67]),
    .in136(pe2neta[68]),
    .in137(pe2netb[68]),
    .in138(pe2neta[69]),
    .in139(pe2netb[69]),
    .in140(pe2neta[70]),
    .in141(pe2netb[70]),
    .in142(pe2neta[71]),
    .in143(pe2netb[71]),
    .in144(pe2neta[72]),
    .in145(pe2netb[72]),
    .in146(pe2neta[73]),
    .in147(pe2netb[73]),
    .in148(pe2neta[74]),
    .in149(pe2netb[74]),
    .in150(pe2neta[75]),
    .in151(pe2netb[75]),
    .in152(pe2neta[76]),
    .in153(pe2netb[76]),
    .in154(pe2neta[77]),
    .in155(pe2netb[77]),
    .in156(pe2neta[78]),
    .in157(pe2netb[78]),
    .in158(pe2neta[79]),
    .in159(pe2netb[79]),
    .in160(pe2neta[80]),
    .in161(pe2netb[80]),
    .in162(pe2neta[81]),
    .in163(pe2netb[81]),
    .in164(pe2neta[82]),
    .in165(pe2netb[82]),
    .in166(pe2neta[83]),
    .in167(pe2netb[83]),
    .in168(pe2neta[84]),
    .in169(pe2netb[84]),
    .in170(pe2neta[85]),
    .in171(pe2netb[85]),
    .in172(pe2neta[86]),
    .in173(pe2netb[86]),
    .in174(pe2neta[87]),
    .in175(pe2netb[87]),
    .in176(pe2neta[88]),
    .in177(pe2netb[88]),
    .in178(pe2neta[89]),
    .in179(pe2netb[89]),
    .in180(pe2neta[90]),
    .in181(pe2netb[90]),
    .in182(pe2neta[91]),
    .in183(pe2netb[91]),
    .in184(pe2neta[92]),
    .in185(pe2netb[92]),
    .in186(pe2neta[93]),
    .in187(pe2netb[93]),
    .in188(pe2neta[94]),
    .in189(pe2netb[94]),
    .in190(pe2neta[95]),
    .in191(pe2netb[95]),
    .in192(pe2neta[96]),
    .in193(pe2netb[96]),
    .in194(pe2neta[97]),
    .in195(pe2netb[97]),
    .in196(pe2neta[98]),
    .in197(pe2netb[98]),
    .in198(pe2neta[99]),
    .in199(pe2netb[99]),
    .in200(pe2neta[100]),
    .in201(pe2netb[100]),
    .in202(pe2neta[101]),
    .in203(pe2netb[101]),
    .in204(pe2neta[102]),
    .in205(pe2netb[102]),
    .in206(pe2neta[103]),
    .in207(pe2netb[103]),
    .in208(pe2neta[104]),
    .in209(pe2netb[104]),
    .in210(pe2neta[105]),
    .in211(pe2netb[105]),
    .in212(pe2neta[106]),
    .in213(pe2netb[106]),
    .in214(pe2neta[107]),
    .in215(pe2netb[107]),
    .in216(pe2neta[108]),
    .in217(pe2netb[108]),
    .in218(pe2neta[109]),
    .in219(pe2netb[109]),
    .in220(pe2neta[110]),
    .in221(pe2netb[110]),
    .in222(pe2neta[111]),
    .in223(pe2netb[111]),
    .in224(pe2neta[112]),
    .in225(pe2netb[112]),
    .in226(pe2neta[113]),
    .in227(pe2netb[113]),
    .in228(pe2neta[114]),
    .in229(pe2netb[114]),
    .in230(pe2neta[115]),
    .in231(pe2netb[115]),
    .in232(pe2neta[116]),
    .in233(pe2netb[116]),
    .in234(pe2neta[117]),
    .in235(pe2netb[117]),
    .in236(pe2neta[118]),
    .in237(pe2netb[118]),
    .in238(pe2neta[119]),
    .in239(pe2netb[119]),
    .in240(pe2neta[120]),
    .in241(pe2netb[120]),
    .in242(pe2neta[121]),
    .in243(pe2netb[121]),
    .in244(pe2neta[122]),
    .in245(pe2netb[122]),
    .in246(pe2neta[123]),
    .in247(pe2netb[123]),
    .in248(pe2neta[124]),
    .in249(pe2netb[124]),
    .in250(pe2neta[125]),
    .in251(pe2netb[125]),
    .in252(pe2neta[126]),
    .in253(pe2netb[126]),
    .in254(pe2neta[127]),
    .in255(pe2netb[127]),
    .out0(net2pea[0]),
    .out1(net2peb[0]),
    .out2(net2pea[1]),
    .out3(net2peb[1]),
    .out4(net2pea[2]),
    .out5(net2peb[2]),
    .out6(net2pea[3]),
    .out7(net2peb[3]),
    .out8(net2pea[4]),
    .out9(net2peb[4]),
    .out10(net2pea[5]),
    .out11(net2peb[5]),
    .out12(net2pea[6]),
    .out13(net2peb[6]),
    .out14(net2pea[7]),
    .out15(net2peb[7]),
    .out16(net2pea[8]),
    .out17(net2peb[8]),
    .out18(net2pea[9]),
    .out19(net2peb[9]),
    .out20(net2pea[10]),
    .out21(net2peb[10]),
    .out22(net2pea[11]),
    .out23(net2peb[11]),
    .out24(net2pea[12]),
    .out25(net2peb[12]),
    .out26(net2pea[13]),
    .out27(net2peb[13]),
    .out28(net2pea[14]),
    .out29(net2peb[14]),
    .out30(net2pea[15]),
    .out31(net2peb[15]),
    .out32(net2pea[16]),
    .out33(net2peb[16]),
    .out34(net2pea[17]),
    .out35(net2peb[17]),
    .out36(net2pea[18]),
    .out37(net2peb[18]),
    .out38(net2pea[19]),
    .out39(net2peb[19]),
    .out40(net2pea[20]),
    .out41(net2peb[20]),
    .out42(net2pea[21]),
    .out43(net2peb[21]),
    .out44(net2pea[22]),
    .out45(net2peb[22]),
    .out46(net2pea[23]),
    .out47(net2peb[23]),
    .out48(net2pea[24]),
    .out49(net2peb[24]),
    .out50(net2pea[25]),
    .out51(net2peb[25]),
    .out52(net2pea[26]),
    .out53(net2peb[26]),
    .out54(net2pea[27]),
    .out55(net2peb[27]),
    .out56(net2pea[28]),
    .out57(net2peb[28]),
    .out58(net2pea[29]),
    .out59(net2peb[29]),
    .out60(net2pea[30]),
    .out61(net2peb[30]),
    .out62(net2pea[31]),
    .out63(net2peb[31]),
    .out64(net2pea[32]),
    .out65(net2peb[32]),
    .out66(net2pea[33]),
    .out67(net2peb[33]),
    .out68(net2pea[34]),
    .out69(net2peb[34]),
    .out70(net2pea[35]),
    .out71(net2peb[35]),
    .out72(net2pea[36]),
    .out73(net2peb[36]),
    .out74(net2pea[37]),
    .out75(net2peb[37]),
    .out76(net2pea[38]),
    .out77(net2peb[38]),
    .out78(net2pea[39]),
    .out79(net2peb[39]),
    .out80(net2pea[40]),
    .out81(net2peb[40]),
    .out82(net2pea[41]),
    .out83(net2peb[41]),
    .out84(net2pea[42]),
    .out85(net2peb[42]),
    .out86(net2pea[43]),
    .out87(net2peb[43]),
    .out88(net2pea[44]),
    .out89(net2peb[44]),
    .out90(net2pea[45]),
    .out91(net2peb[45]),
    .out92(net2pea[46]),
    .out93(net2peb[46]),
    .out94(net2pea[47]),
    .out95(net2peb[47]),
    .out96(net2pea[48]),
    .out97(net2peb[48]),
    .out98(net2pea[49]),
    .out99(net2peb[49]),
    .out100(net2pea[50]),
    .out101(net2peb[50]),
    .out102(net2pea[51]),
    .out103(net2peb[51]),
    .out104(net2pea[52]),
    .out105(net2peb[52]),
    .out106(net2pea[53]),
    .out107(net2peb[53]),
    .out108(net2pea[54]),
    .out109(net2peb[54]),
    .out110(net2pea[55]),
    .out111(net2peb[55]),
    .out112(net2pea[56]),
    .out113(net2peb[56]),
    .out114(net2pea[57]),
    .out115(net2peb[57]),
    .out116(net2pea[58]),
    .out117(net2peb[58]),
    .out118(net2pea[59]),
    .out119(net2peb[59]),
    .out120(net2pea[60]),
    .out121(net2peb[60]),
    .out122(net2pea[61]),
    .out123(net2peb[61]),
    .out124(net2pea[62]),
    .out125(net2peb[62]),
    .out126(net2pea[63]),
    .out127(net2peb[63]),
    .out128(net2pea[64]),
    .out129(net2peb[64]),
    .out130(net2pea[65]),
    .out131(net2peb[65]),
    .out132(net2pea[66]),
    .out133(net2peb[66]),
    .out134(net2pea[67]),
    .out135(net2peb[67]),
    .out136(net2pea[68]),
    .out137(net2peb[68]),
    .out138(net2pea[69]),
    .out139(net2peb[69]),
    .out140(net2pea[70]),
    .out141(net2peb[70]),
    .out142(net2pea[71]),
    .out143(net2peb[71]),
    .out144(net2pea[72]),
    .out145(net2peb[72]),
    .out146(net2pea[73]),
    .out147(net2peb[73]),
    .out148(net2pea[74]),
    .out149(net2peb[74]),
    .out150(net2pea[75]),
    .out151(net2peb[75]),
    .out152(net2pea[76]),
    .out153(net2peb[76]),
    .out154(net2pea[77]),
    .out155(net2peb[77]),
    .out156(net2pea[78]),
    .out157(net2peb[78]),
    .out158(net2pea[79]),
    .out159(net2peb[79]),
    .out160(net2pea[80]),
    .out161(net2peb[80]),
    .out162(net2pea[81]),
    .out163(net2peb[81]),
    .out164(net2pea[82]),
    .out165(net2peb[82]),
    .out166(net2pea[83]),
    .out167(net2peb[83]),
    .out168(net2pea[84]),
    .out169(net2peb[84]),
    .out170(net2pea[85]),
    .out171(net2peb[85]),
    .out172(net2pea[86]),
    .out173(net2peb[86]),
    .out174(net2pea[87]),
    .out175(net2peb[87]),
    .out176(net2pea[88]),
    .out177(net2peb[88]),
    .out178(net2pea[89]),
    .out179(net2peb[89]),
    .out180(net2pea[90]),
    .out181(net2peb[90]),
    .out182(net2pea[91]),
    .out183(net2peb[91]),
    .out184(net2pea[92]),
    .out185(net2peb[92]),
    .out186(net2pea[93]),
    .out187(net2peb[93]),
    .out188(net2pea[94]),
    .out189(net2peb[94]),
    .out190(net2pea[95]),
    .out191(net2peb[95]),
    .out192(net2pea[96]),
    .out193(net2peb[96]),
    .out194(net2pea[97]),
    .out195(net2peb[97]),
    .out196(net2pea[98]),
    .out197(net2peb[98]),
    .out198(net2pea[99]),
    .out199(net2peb[99]),
    .out200(net2pea[100]),
    .out201(net2peb[100]),
    .out202(net2pea[101]),
    .out203(net2peb[101]),
    .out204(net2pea[102]),
    .out205(net2peb[102]),
    .out206(net2pea[103]),
    .out207(net2peb[103]),
    .out208(net2pea[104]),
    .out209(net2peb[104]),
    .out210(net2pea[105]),
    .out211(net2peb[105]),
    .out212(net2pea[106]),
    .out213(net2peb[106]),
    .out214(net2pea[107]),
    .out215(net2peb[107]),
    .out216(net2pea[108]),
    .out217(net2peb[108]),
    .out218(net2pea[109]),
    .out219(net2peb[109]),
    .out220(net2pea[110]),
    .out221(net2peb[110]),
    .out222(net2pea[111]),
    .out223(net2peb[111]),
    .out224(net2pea[112]),
    .out225(net2peb[112]),
    .out226(net2pea[113]),
    .out227(net2peb[113]),
    .out228(net2pea[114]),
    .out229(net2peb[114]),
    .out230(net2pea[115]),
    .out231(net2peb[115]),
    .out232(net2pea[116]),
    .out233(net2peb[116]),
    .out234(net2pea[117]),
    .out235(net2peb[117]),
    .out236(net2pea[118]),
    .out237(net2peb[118]),
    .out238(net2pea[119]),
    .out239(net2peb[119]),
    .out240(net2pea[120]),
    .out241(net2peb[120]),
    .out242(net2pea[121]),
    .out243(net2peb[121]),
    .out244(net2pea[122]),
    .out245(net2peb[122]),
    .out246(net2pea[123]),
    .out247(net2peb[123]),
    .out248(net2pea[124]),
    .out249(net2peb[124]),
    .out250(net2pea[125]),
    .out251(net2peb[125]),
    .out252(net2pea[126]),
    .out253(net2peb[126]),
    .out254(net2pea[127]),
    .out255(net2peb[127])
  );

endmodule