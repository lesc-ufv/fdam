module fir1632(
  input clk,
  input rst,
  input start,
  input [32-1:0] num_conf,
  input [32-1:0] num_data_in,
  input [32-1:0] num_data_out,
  input available_write,
  input available_read,
  output req_rd_data,
  input [512-1:0] rd_data,
  output req_wr_data,
  output [512-1:0] wr_data,
  output done
  );

 wire rdy, en;
 wire [31:0] dconf;
 wire rin1,rin2,rin3,rin4,rin5,rin6,rin7,rin8,rin9,rin10,rin11,rin12,rin13,rin14,rin15,rin16,rin17,rin18,rin19,rin20,rin21,rin22,rin23,rin24,rin25,rin26,rin27,rin28,rin29,rin30,rin31,rin32;
 wire rout1,rout2,rout3,rout4,rout5,rout6,rout7,rout8,rout9,rout10,rout11,rout12,rout13,rout14,rout15,rout16,rout17,rout18,rout19,rout20,rout21,rout22,rout23,rout24,rout25,rout26,rout27,rout28,rout29,rout30,rout31,rout32;
 wire [15:0] din1,din2,din3,din4,din5,din6,din7,din8,din9,din10,din11,din12,din13,din14,din15,din16,din17,din18,din19,din20,din21,din22,din23,din24,din25,din26,din27,din28,din29,din30,din31,din32;
 wire [15:0] dout1,dout2,dout3,dout4,dout5,dout6,dout7,dout8,dout9,dout10,dout11,dout12,dout13,dout14,dout15,dout16,dout17,dout18,dout19,dout20,dout21,dout22,dout23,dout24,dout25,dout26,dout27,dout28,dout29,dout30,dout31,dout32;
  
hebe_in32
hebe_in32_
(
  .clk(clk),
  .rst(rst),
  .start(start),
  .num_data(num_data_in),
  .num_conf(num_conf),
  .rdy(rdy),
  .available_read(available_read),
  .rd_data(rd_data),
  .req_rd_data(req_rd_data),
  .dconf(dconf),
  .en(en),
  .rout1(rin1),
  .rout2(rin2),
  .rout3(rin3),
  .rout4(rin4),
  .rout5(rin5),
  .rout6(rin6),
  .rout7(rin7),
  .rout8(rin8),
  .rout9(rin9),
  .rout10(rin10),
  .rout11(rin11),
  .rout12(rin12),
  .rout13(rin13),
  .rout14(rin14),
  .rout15(rin15),
  .rout16(rin16),
  .rout17(rin17),
  .rout18(rin18),
  .rout19(rin19),
  .rout20(rin20),
  .rout21(rin21),
  .rout22(rin22),
  .rout23(rin23),
  .rout24(rin24),
  .rout25(rin25),
  .rout26(rin26),
  .rout27(rin27),
  .rout28(rin28),
  .rout29(rin29),
  .rout30(rin30),
  .rout31(rin31),
  .rout32(rin32),
  .dout1(din1),
  .dout2(din2),
  .dout3(din3),
  .dout4(din4),
  .dout5(din5),
  .dout6(din6),
  .dout7(din7),
  .dout8(din8),
  .dout9(din9),
  .dout10(din10),
  .dout11(din11),
  .dout12(din12),
  .dout13(din13),
  .dout14(din14),
  .dout15(din15),
  .dout16(din16),
  .dout17(din17),
  .dout18(din18),
  .dout19(din19),
  .dout20(din20),
  .dout21(din21),
  .dout22(din22),
  .dout23(din23),
  .dout24(din24),
  .dout25(din25),
  .dout26(din26),
  .dout27(din27),
  .dout28(din28),
  .dout29(din29),
  .dout30(din30),
  .dout31(din31),
  .dout32(din32)
);
  

hebe_out32
hebe_out32_
(
  .clk(clk),
  .rst(rst),
  .start(start),
  .num_data(num_data_out),
  .en(en),
  .rin1(rout1),
  .rin2(rout2),
  .rin3(rout3),
  .rin4(rout4),
  .rin5(rout5),
  .rin6(rout6),
  .rin7(rout7),
  .rin8(rout8),
  .rin9(rout9),
  .rin10(rout10),
  .rin11(rout11),
  .rin12(rout12),
  .rin13(rout13),
  .rin14(rout14),
  .rin15(rout15),
  .rin16(rout16),
  .rin17(rout17),
  .rin18(rout18),
  .rin19(rout19),
  .rin20(rout20),
  .rin21(rout21),
  .rin22(rout22),
  .rin23(rout23),
  .rin24(rout24),
  .rin25(rout25),
  .rin26(rout26),
  .rin27(rout27),
  .rin28(rout28),
  .rin29(rout29),
  .rin30(rout30),
  .rin31(rout31),
  .rin32(rout32),
  .din1(dout1),
  .din2(dout2),
  .din3(dout3),
  .din4(dout4),
  .din5(dout5),
  .din6(dout6),
  .din7(dout7),
  .din8(dout8),
  .din9(dout9),
  .din10(dout10),
  .din11(dout11),
  .din12(dout12),
  .din13(dout13),
  .din14(dout14),
  .din15(dout15),
  .din16(dout16),
  .din17(dout17),
  .din18(dout18),
  .din19(dout19),
  .din20(dout20),
  .din21(dout21),
  .din22(dout22),
  .din23(dout23),
  .din24(dout24),
  .din25(dout25),
  .din26(dout26),
  .din27(dout27),
  .din28(dout28),
  .din29(dout29),
  .din30(dout30),
  .din31(dout31),
  .din32(dout32),
  .available_write(available_write),
  .req_wr_data(req_wr_data),
  .wr_data(wr_data),
  .rdy(rdy),
  .done(done)
);  
  

fir16
fir16_1
(
  .clk(clk),
  .rst(rst),
  .din(din1),
  .rin(rin1),
  .dconf(dconf),
  .dout(dout1),
  .rout(rout1),
  .en(en)
);

fir16
fir16_2
(
  .clk(clk),
  .rst(rst),
  .din(din2),
  .rin(rin2),
  .dconf(dconf),
  .dout(dout2),
  .rout(rout2),
  .en(en)
);

fir16
fir16_3
(
  .clk(clk),
  .rst(rst),
  .din(din3),
  .rin(rin3),
  .dconf(dconf),
  .dout(dout3),
  .rout(rout3),
  .en(en)
);

fir16
fir16_4
(
  .clk(clk),
  .rst(rst),
  .din(din4),
  .rin(rin4),
  .dconf(dconf),
  .dout(dout4),
  .rout(rout4),
  .en(en)
);

fir16
fir16_5
(
  .clk(clk),
  .rst(rst),
  .din(din5),
  .rin(rin5),
  .dconf(dconf),
  .dout(dout5),
  .rout(rout5),
  .en(en)
);

fir16
fir16_6
(
  .clk(clk),
  .rst(rst),
  .din(din6),
  .rin(rin6),
  .dconf(dconf),
  .dout(dout6),
  .rout(rout6),
  .en(en)
);

fir16
fir16_7
(
  .clk(clk),
  .rst(rst),
  .din(din7),
  .rin(rin7),
  .dconf(dconf),
  .dout(dout7),
  .rout(rout7),
  .en(en)
);

fir16
fir16_8
(
  .clk(clk),
  .rst(rst),
  .din(din8),
  .rin(rin8),
  .dconf(dconf),
  .dout(dout8),
  .rout(rout8),
  .en(en)
);

fir16
fir16_9
(
  .clk(clk),
  .rst(rst),
  .din(din9),
  .rin(rin9),
  .dconf(dconf),
  .dout(dout9),
  .rout(rout9),
  .en(en)
);

fir16
fir16_10
(
  .clk(clk),
  .rst(rst),
  .din(din10),
  .rin(rin10),
  .dconf(dconf),
  .dout(dout10),
  .rout(rout10),
  .en(en)
);

fir16
fir16_11
(
  .clk(clk),
  .rst(rst),
  .din(din11),
  .rin(rin11),
  .dconf(dconf),
  .dout(dout11),
  .rout(rout11),
  .en(en)
);

fir16
fir16_12
(
  .clk(clk),
  .rst(rst),
  .din(din12),
  .rin(rin12),
  .dconf(dconf),
  .dout(dout12),
  .rout(rout12),
  .en(en)
);

fir16
fir16_13
(
  .clk(clk),
  .rst(rst),
  .din(din13),
  .rin(rin13),
  .dconf(dconf),
  .dout(dout13),
  .rout(rout13),
  .en(en)
);

fir16
fir16_14
(
  .clk(clk),
  .rst(rst),
  .din(din14),
  .rin(rin14),
  .dconf(dconf),
  .dout(dout14),
  .rout(rout14),
  .en(en)
);

fir16
fir16_15
(
  .clk(clk),
  .rst(rst),
  .din(din15),
  .rin(rin15),
  .dconf(dconf),
  .dout(dout15),
  .rout(rout15),
  .en(en)
);

fir16
fir16_16
(
  .clk(clk),
  .rst(rst),
  .din(din16),
  .rin(rin16),
  .dconf(dconf),
  .dout(dout16),
  .rout(rout16),
  .en(en)
);

fir16
fir16_17
(
  .clk(clk),
  .rst(rst),
  .din(din17),
  .rin(rin17),
  .dconf(dconf),
  .dout(dout17),
  .rout(rout17),
  .en(en)
);

fir16
fir16_18
(
  .clk(clk),
  .rst(rst),
  .din(din18),
  .rin(rin18),
  .dconf(dconf),
  .dout(dout18),
  .rout(rout18),
  .en(en)
);

fir16
fir16_19
(
  .clk(clk),
  .rst(rst),
  .din(din19),
  .rin(rin19),
  .dconf(dconf),
  .dout(dout19),
  .rout(rout19),
  .en(en)
);

fir16
fir16_20
(
  .clk(clk),
  .rst(rst),
  .din(din20),
  .rin(rin20),
  .dconf(dconf),
  .dout(dout20),
  .rout(rout20),
  .en(en)
);

fir16
fir16_21
(
  .clk(clk),
  .rst(rst),
  .din(din21),
  .rin(rin21),
  .dconf(dconf),
  .dout(dout21),
  .rout(rout21),
  .en(en)
);

fir16
fir16_22
(
  .clk(clk),
  .rst(rst),
  .din(din22),
  .rin(rin22),
  .dconf(dconf),
  .dout(dout22),
  .rout(rout22),
  .en(en)
);

fir16
fir16_23
(
  .clk(clk),
  .rst(rst),
  .din(din23),
  .rin(rin23),
  .dconf(dconf),
  .dout(dout23),
  .rout(rout23),
  .en(en)
);

fir16
fir16_24
(
  .clk(clk),
  .rst(rst),
  .din(din24),
  .rin(rin24),
  .dconf(dconf),
  .dout(dout24),
  .rout(rout24),
  .en(en)
);

fir16
fir16_25
(
  .clk(clk),
  .rst(rst),
  .din(din25),
  .rin(rin25),
  .dconf(dconf),
  .dout(dout25),
  .rout(rout25),
  .en(en)
);

fir16
fir16_26
(
  .clk(clk),
  .rst(rst),
  .din(din26),
  .rin(rin26),
  .dconf(dconf),
  .dout(dout26),
  .rout(rout26),
  .en(en)
);

fir16
fir16_27
(
  .clk(clk),
  .rst(rst),
  .din(din27),
  .rin(rin27),
  .dconf(dconf),
  .dout(dout27),
  .rout(rout27),
  .en(en)
);

fir16
fir16_28
(
  .clk(clk),
  .rst(rst),
  .din(din28),
  .rin(rin28),
  .dconf(dconf),
  .dout(dout28),
  .rout(rout28),
  .en(en)
);

fir16
fir16_29
(
  .clk(clk),
  .rst(rst),
  .din(din29),
  .rin(rin29),
  .dconf(dconf),
  .dout(dout29),
  .rout(rout29),
  .en(en)
);

fir16
fir16_30
(
  .clk(clk),
  .rst(rst),
  .din(din30),
  .rin(rin30),
  .dconf(dconf),
  .dout(dout30),
  .rout(rout30),
  .en(en)
);

fir16
fir16_31
(
  .clk(clk),
  .rst(rst),
  .din(din31),
  .rin(rin31),
  .dconf(dconf),
  .dout(dout31),
  .rout(rout31),
  .en(en)
);

fir16
fir16_32
(
  .clk(clk),
  .rst(rst),
  .din(din32),
  .rin(rin32),
  .dconf(dconf),
  .dout(dout32),
  .rout(rout32),
  .en(en)
);

endmodule
