module omega256x256_4_0_8 #
(
  parameter WIDTH = 16,
  parameter PIPE_EXTRA = 0
)
(
  input clk,
  input rst,
  input [256-1:0] en_pc_net,
  input [1280-1:0] en,
  input [64-1:0] net_conf_bus_in,
  input [WIDTH-1:0] in0,
  input [WIDTH-1:0] in1,
  input [WIDTH-1:0] in2,
  input [WIDTH-1:0] in3,
  input [WIDTH-1:0] in4,
  input [WIDTH-1:0] in5,
  input [WIDTH-1:0] in6,
  input [WIDTH-1:0] in7,
  input [WIDTH-1:0] in8,
  input [WIDTH-1:0] in9,
  input [WIDTH-1:0] in10,
  input [WIDTH-1:0] in11,
  input [WIDTH-1:0] in12,
  input [WIDTH-1:0] in13,
  input [WIDTH-1:0] in14,
  input [WIDTH-1:0] in15,
  input [WIDTH-1:0] in16,
  input [WIDTH-1:0] in17,
  input [WIDTH-1:0] in18,
  input [WIDTH-1:0] in19,
  input [WIDTH-1:0] in20,
  input [WIDTH-1:0] in21,
  input [WIDTH-1:0] in22,
  input [WIDTH-1:0] in23,
  input [WIDTH-1:0] in24,
  input [WIDTH-1:0] in25,
  input [WIDTH-1:0] in26,
  input [WIDTH-1:0] in27,
  input [WIDTH-1:0] in28,
  input [WIDTH-1:0] in29,
  input [WIDTH-1:0] in30,
  input [WIDTH-1:0] in31,
  input [WIDTH-1:0] in32,
  input [WIDTH-1:0] in33,
  input [WIDTH-1:0] in34,
  input [WIDTH-1:0] in35,
  input [WIDTH-1:0] in36,
  input [WIDTH-1:0] in37,
  input [WIDTH-1:0] in38,
  input [WIDTH-1:0] in39,
  input [WIDTH-1:0] in40,
  input [WIDTH-1:0] in41,
  input [WIDTH-1:0] in42,
  input [WIDTH-1:0] in43,
  input [WIDTH-1:0] in44,
  input [WIDTH-1:0] in45,
  input [WIDTH-1:0] in46,
  input [WIDTH-1:0] in47,
  input [WIDTH-1:0] in48,
  input [WIDTH-1:0] in49,
  input [WIDTH-1:0] in50,
  input [WIDTH-1:0] in51,
  input [WIDTH-1:0] in52,
  input [WIDTH-1:0] in53,
  input [WIDTH-1:0] in54,
  input [WIDTH-1:0] in55,
  input [WIDTH-1:0] in56,
  input [WIDTH-1:0] in57,
  input [WIDTH-1:0] in58,
  input [WIDTH-1:0] in59,
  input [WIDTH-1:0] in60,
  input [WIDTH-1:0] in61,
  input [WIDTH-1:0] in62,
  input [WIDTH-1:0] in63,
  input [WIDTH-1:0] in64,
  input [WIDTH-1:0] in65,
  input [WIDTH-1:0] in66,
  input [WIDTH-1:0] in67,
  input [WIDTH-1:0] in68,
  input [WIDTH-1:0] in69,
  input [WIDTH-1:0] in70,
  input [WIDTH-1:0] in71,
  input [WIDTH-1:0] in72,
  input [WIDTH-1:0] in73,
  input [WIDTH-1:0] in74,
  input [WIDTH-1:0] in75,
  input [WIDTH-1:0] in76,
  input [WIDTH-1:0] in77,
  input [WIDTH-1:0] in78,
  input [WIDTH-1:0] in79,
  input [WIDTH-1:0] in80,
  input [WIDTH-1:0] in81,
  input [WIDTH-1:0] in82,
  input [WIDTH-1:0] in83,
  input [WIDTH-1:0] in84,
  input [WIDTH-1:0] in85,
  input [WIDTH-1:0] in86,
  input [WIDTH-1:0] in87,
  input [WIDTH-1:0] in88,
  input [WIDTH-1:0] in89,
  input [WIDTH-1:0] in90,
  input [WIDTH-1:0] in91,
  input [WIDTH-1:0] in92,
  input [WIDTH-1:0] in93,
  input [WIDTH-1:0] in94,
  input [WIDTH-1:0] in95,
  input [WIDTH-1:0] in96,
  input [WIDTH-1:0] in97,
  input [WIDTH-1:0] in98,
  input [WIDTH-1:0] in99,
  input [WIDTH-1:0] in100,
  input [WIDTH-1:0] in101,
  input [WIDTH-1:0] in102,
  input [WIDTH-1:0] in103,
  input [WIDTH-1:0] in104,
  input [WIDTH-1:0] in105,
  input [WIDTH-1:0] in106,
  input [WIDTH-1:0] in107,
  input [WIDTH-1:0] in108,
  input [WIDTH-1:0] in109,
  input [WIDTH-1:0] in110,
  input [WIDTH-1:0] in111,
  input [WIDTH-1:0] in112,
  input [WIDTH-1:0] in113,
  input [WIDTH-1:0] in114,
  input [WIDTH-1:0] in115,
  input [WIDTH-1:0] in116,
  input [WIDTH-1:0] in117,
  input [WIDTH-1:0] in118,
  input [WIDTH-1:0] in119,
  input [WIDTH-1:0] in120,
  input [WIDTH-1:0] in121,
  input [WIDTH-1:0] in122,
  input [WIDTH-1:0] in123,
  input [WIDTH-1:0] in124,
  input [WIDTH-1:0] in125,
  input [WIDTH-1:0] in126,
  input [WIDTH-1:0] in127,
  input [WIDTH-1:0] in128,
  input [WIDTH-1:0] in129,
  input [WIDTH-1:0] in130,
  input [WIDTH-1:0] in131,
  input [WIDTH-1:0] in132,
  input [WIDTH-1:0] in133,
  input [WIDTH-1:0] in134,
  input [WIDTH-1:0] in135,
  input [WIDTH-1:0] in136,
  input [WIDTH-1:0] in137,
  input [WIDTH-1:0] in138,
  input [WIDTH-1:0] in139,
  input [WIDTH-1:0] in140,
  input [WIDTH-1:0] in141,
  input [WIDTH-1:0] in142,
  input [WIDTH-1:0] in143,
  input [WIDTH-1:0] in144,
  input [WIDTH-1:0] in145,
  input [WIDTH-1:0] in146,
  input [WIDTH-1:0] in147,
  input [WIDTH-1:0] in148,
  input [WIDTH-1:0] in149,
  input [WIDTH-1:0] in150,
  input [WIDTH-1:0] in151,
  input [WIDTH-1:0] in152,
  input [WIDTH-1:0] in153,
  input [WIDTH-1:0] in154,
  input [WIDTH-1:0] in155,
  input [WIDTH-1:0] in156,
  input [WIDTH-1:0] in157,
  input [WIDTH-1:0] in158,
  input [WIDTH-1:0] in159,
  input [WIDTH-1:0] in160,
  input [WIDTH-1:0] in161,
  input [WIDTH-1:0] in162,
  input [WIDTH-1:0] in163,
  input [WIDTH-1:0] in164,
  input [WIDTH-1:0] in165,
  input [WIDTH-1:0] in166,
  input [WIDTH-1:0] in167,
  input [WIDTH-1:0] in168,
  input [WIDTH-1:0] in169,
  input [WIDTH-1:0] in170,
  input [WIDTH-1:0] in171,
  input [WIDTH-1:0] in172,
  input [WIDTH-1:0] in173,
  input [WIDTH-1:0] in174,
  input [WIDTH-1:0] in175,
  input [WIDTH-1:0] in176,
  input [WIDTH-1:0] in177,
  input [WIDTH-1:0] in178,
  input [WIDTH-1:0] in179,
  input [WIDTH-1:0] in180,
  input [WIDTH-1:0] in181,
  input [WIDTH-1:0] in182,
  input [WIDTH-1:0] in183,
  input [WIDTH-1:0] in184,
  input [WIDTH-1:0] in185,
  input [WIDTH-1:0] in186,
  input [WIDTH-1:0] in187,
  input [WIDTH-1:0] in188,
  input [WIDTH-1:0] in189,
  input [WIDTH-1:0] in190,
  input [WIDTH-1:0] in191,
  input [WIDTH-1:0] in192,
  input [WIDTH-1:0] in193,
  input [WIDTH-1:0] in194,
  input [WIDTH-1:0] in195,
  input [WIDTH-1:0] in196,
  input [WIDTH-1:0] in197,
  input [WIDTH-1:0] in198,
  input [WIDTH-1:0] in199,
  input [WIDTH-1:0] in200,
  input [WIDTH-1:0] in201,
  input [WIDTH-1:0] in202,
  input [WIDTH-1:0] in203,
  input [WIDTH-1:0] in204,
  input [WIDTH-1:0] in205,
  input [WIDTH-1:0] in206,
  input [WIDTH-1:0] in207,
  input [WIDTH-1:0] in208,
  input [WIDTH-1:0] in209,
  input [WIDTH-1:0] in210,
  input [WIDTH-1:0] in211,
  input [WIDTH-1:0] in212,
  input [WIDTH-1:0] in213,
  input [WIDTH-1:0] in214,
  input [WIDTH-1:0] in215,
  input [WIDTH-1:0] in216,
  input [WIDTH-1:0] in217,
  input [WIDTH-1:0] in218,
  input [WIDTH-1:0] in219,
  input [WIDTH-1:0] in220,
  input [WIDTH-1:0] in221,
  input [WIDTH-1:0] in222,
  input [WIDTH-1:0] in223,
  input [WIDTH-1:0] in224,
  input [WIDTH-1:0] in225,
  input [WIDTH-1:0] in226,
  input [WIDTH-1:0] in227,
  input [WIDTH-1:0] in228,
  input [WIDTH-1:0] in229,
  input [WIDTH-1:0] in230,
  input [WIDTH-1:0] in231,
  input [WIDTH-1:0] in232,
  input [WIDTH-1:0] in233,
  input [WIDTH-1:0] in234,
  input [WIDTH-1:0] in235,
  input [WIDTH-1:0] in236,
  input [WIDTH-1:0] in237,
  input [WIDTH-1:0] in238,
  input [WIDTH-1:0] in239,
  input [WIDTH-1:0] in240,
  input [WIDTH-1:0] in241,
  input [WIDTH-1:0] in242,
  input [WIDTH-1:0] in243,
  input [WIDTH-1:0] in244,
  input [WIDTH-1:0] in245,
  input [WIDTH-1:0] in246,
  input [WIDTH-1:0] in247,
  input [WIDTH-1:0] in248,
  input [WIDTH-1:0] in249,
  input [WIDTH-1:0] in250,
  input [WIDTH-1:0] in251,
  input [WIDTH-1:0] in252,
  input [WIDTH-1:0] in253,
  input [WIDTH-1:0] in254,
  input [WIDTH-1:0] in255,
  output [WIDTH-1:0] out0,
  output [WIDTH-1:0] out1,
  output [WIDTH-1:0] out2,
  output [WIDTH-1:0] out3,
  output [WIDTH-1:0] out4,
  output [WIDTH-1:0] out5,
  output [WIDTH-1:0] out6,
  output [WIDTH-1:0] out7,
  output [WIDTH-1:0] out8,
  output [WIDTH-1:0] out9,
  output [WIDTH-1:0] out10,
  output [WIDTH-1:0] out11,
  output [WIDTH-1:0] out12,
  output [WIDTH-1:0] out13,
  output [WIDTH-1:0] out14,
  output [WIDTH-1:0] out15,
  output [WIDTH-1:0] out16,
  output [WIDTH-1:0] out17,
  output [WIDTH-1:0] out18,
  output [WIDTH-1:0] out19,
  output [WIDTH-1:0] out20,
  output [WIDTH-1:0] out21,
  output [WIDTH-1:0] out22,
  output [WIDTH-1:0] out23,
  output [WIDTH-1:0] out24,
  output [WIDTH-1:0] out25,
  output [WIDTH-1:0] out26,
  output [WIDTH-1:0] out27,
  output [WIDTH-1:0] out28,
  output [WIDTH-1:0] out29,
  output [WIDTH-1:0] out30,
  output [WIDTH-1:0] out31,
  output [WIDTH-1:0] out32,
  output [WIDTH-1:0] out33,
  output [WIDTH-1:0] out34,
  output [WIDTH-1:0] out35,
  output [WIDTH-1:0] out36,
  output [WIDTH-1:0] out37,
  output [WIDTH-1:0] out38,
  output [WIDTH-1:0] out39,
  output [WIDTH-1:0] out40,
  output [WIDTH-1:0] out41,
  output [WIDTH-1:0] out42,
  output [WIDTH-1:0] out43,
  output [WIDTH-1:0] out44,
  output [WIDTH-1:0] out45,
  output [WIDTH-1:0] out46,
  output [WIDTH-1:0] out47,
  output [WIDTH-1:0] out48,
  output [WIDTH-1:0] out49,
  output [WIDTH-1:0] out50,
  output [WIDTH-1:0] out51,
  output [WIDTH-1:0] out52,
  output [WIDTH-1:0] out53,
  output [WIDTH-1:0] out54,
  output [WIDTH-1:0] out55,
  output [WIDTH-1:0] out56,
  output [WIDTH-1:0] out57,
  output [WIDTH-1:0] out58,
  output [WIDTH-1:0] out59,
  output [WIDTH-1:0] out60,
  output [WIDTH-1:0] out61,
  output [WIDTH-1:0] out62,
  output [WIDTH-1:0] out63,
  output [WIDTH-1:0] out64,
  output [WIDTH-1:0] out65,
  output [WIDTH-1:0] out66,
  output [WIDTH-1:0] out67,
  output [WIDTH-1:0] out68,
  output [WIDTH-1:0] out69,
  output [WIDTH-1:0] out70,
  output [WIDTH-1:0] out71,
  output [WIDTH-1:0] out72,
  output [WIDTH-1:0] out73,
  output [WIDTH-1:0] out74,
  output [WIDTH-1:0] out75,
  output [WIDTH-1:0] out76,
  output [WIDTH-1:0] out77,
  output [WIDTH-1:0] out78,
  output [WIDTH-1:0] out79,
  output [WIDTH-1:0] out80,
  output [WIDTH-1:0] out81,
  output [WIDTH-1:0] out82,
  output [WIDTH-1:0] out83,
  output [WIDTH-1:0] out84,
  output [WIDTH-1:0] out85,
  output [WIDTH-1:0] out86,
  output [WIDTH-1:0] out87,
  output [WIDTH-1:0] out88,
  output [WIDTH-1:0] out89,
  output [WIDTH-1:0] out90,
  output [WIDTH-1:0] out91,
  output [WIDTH-1:0] out92,
  output [WIDTH-1:0] out93,
  output [WIDTH-1:0] out94,
  output [WIDTH-1:0] out95,
  output [WIDTH-1:0] out96,
  output [WIDTH-1:0] out97,
  output [WIDTH-1:0] out98,
  output [WIDTH-1:0] out99,
  output [WIDTH-1:0] out100,
  output [WIDTH-1:0] out101,
  output [WIDTH-1:0] out102,
  output [WIDTH-1:0] out103,
  output [WIDTH-1:0] out104,
  output [WIDTH-1:0] out105,
  output [WIDTH-1:0] out106,
  output [WIDTH-1:0] out107,
  output [WIDTH-1:0] out108,
  output [WIDTH-1:0] out109,
  output [WIDTH-1:0] out110,
  output [WIDTH-1:0] out111,
  output [WIDTH-1:0] out112,
  output [WIDTH-1:0] out113,
  output [WIDTH-1:0] out114,
  output [WIDTH-1:0] out115,
  output [WIDTH-1:0] out116,
  output [WIDTH-1:0] out117,
  output [WIDTH-1:0] out118,
  output [WIDTH-1:0] out119,
  output [WIDTH-1:0] out120,
  output [WIDTH-1:0] out121,
  output [WIDTH-1:0] out122,
  output [WIDTH-1:0] out123,
  output [WIDTH-1:0] out124,
  output [WIDTH-1:0] out125,
  output [WIDTH-1:0] out126,
  output [WIDTH-1:0] out127,
  output [WIDTH-1:0] out128,
  output [WIDTH-1:0] out129,
  output [WIDTH-1:0] out130,
  output [WIDTH-1:0] out131,
  output [WIDTH-1:0] out132,
  output [WIDTH-1:0] out133,
  output [WIDTH-1:0] out134,
  output [WIDTH-1:0] out135,
  output [WIDTH-1:0] out136,
  output [WIDTH-1:0] out137,
  output [WIDTH-1:0] out138,
  output [WIDTH-1:0] out139,
  output [WIDTH-1:0] out140,
  output [WIDTH-1:0] out141,
  output [WIDTH-1:0] out142,
  output [WIDTH-1:0] out143,
  output [WIDTH-1:0] out144,
  output [WIDTH-1:0] out145,
  output [WIDTH-1:0] out146,
  output [WIDTH-1:0] out147,
  output [WIDTH-1:0] out148,
  output [WIDTH-1:0] out149,
  output [WIDTH-1:0] out150,
  output [WIDTH-1:0] out151,
  output [WIDTH-1:0] out152,
  output [WIDTH-1:0] out153,
  output [WIDTH-1:0] out154,
  output [WIDTH-1:0] out155,
  output [WIDTH-1:0] out156,
  output [WIDTH-1:0] out157,
  output [WIDTH-1:0] out158,
  output [WIDTH-1:0] out159,
  output [WIDTH-1:0] out160,
  output [WIDTH-1:0] out161,
  output [WIDTH-1:0] out162,
  output [WIDTH-1:0] out163,
  output [WIDTH-1:0] out164,
  output [WIDTH-1:0] out165,
  output [WIDTH-1:0] out166,
  output [WIDTH-1:0] out167,
  output [WIDTH-1:0] out168,
  output [WIDTH-1:0] out169,
  output [WIDTH-1:0] out170,
  output [WIDTH-1:0] out171,
  output [WIDTH-1:0] out172,
  output [WIDTH-1:0] out173,
  output [WIDTH-1:0] out174,
  output [WIDTH-1:0] out175,
  output [WIDTH-1:0] out176,
  output [WIDTH-1:0] out177,
  output [WIDTH-1:0] out178,
  output [WIDTH-1:0] out179,
  output [WIDTH-1:0] out180,
  output [WIDTH-1:0] out181,
  output [WIDTH-1:0] out182,
  output [WIDTH-1:0] out183,
  output [WIDTH-1:0] out184,
  output [WIDTH-1:0] out185,
  output [WIDTH-1:0] out186,
  output [WIDTH-1:0] out187,
  output [WIDTH-1:0] out188,
  output [WIDTH-1:0] out189,
  output [WIDTH-1:0] out190,
  output [WIDTH-1:0] out191,
  output [WIDTH-1:0] out192,
  output [WIDTH-1:0] out193,
  output [WIDTH-1:0] out194,
  output [WIDTH-1:0] out195,
  output [WIDTH-1:0] out196,
  output [WIDTH-1:0] out197,
  output [WIDTH-1:0] out198,
  output [WIDTH-1:0] out199,
  output [WIDTH-1:0] out200,
  output [WIDTH-1:0] out201,
  output [WIDTH-1:0] out202,
  output [WIDTH-1:0] out203,
  output [WIDTH-1:0] out204,
  output [WIDTH-1:0] out205,
  output [WIDTH-1:0] out206,
  output [WIDTH-1:0] out207,
  output [WIDTH-1:0] out208,
  output [WIDTH-1:0] out209,
  output [WIDTH-1:0] out210,
  output [WIDTH-1:0] out211,
  output [WIDTH-1:0] out212,
  output [WIDTH-1:0] out213,
  output [WIDTH-1:0] out214,
  output [WIDTH-1:0] out215,
  output [WIDTH-1:0] out216,
  output [WIDTH-1:0] out217,
  output [WIDTH-1:0] out218,
  output [WIDTH-1:0] out219,
  output [WIDTH-1:0] out220,
  output [WIDTH-1:0] out221,
  output [WIDTH-1:0] out222,
  output [WIDTH-1:0] out223,
  output [WIDTH-1:0] out224,
  output [WIDTH-1:0] out225,
  output [WIDTH-1:0] out226,
  output [WIDTH-1:0] out227,
  output [WIDTH-1:0] out228,
  output [WIDTH-1:0] out229,
  output [WIDTH-1:0] out230,
  output [WIDTH-1:0] out231,
  output [WIDTH-1:0] out232,
  output [WIDTH-1:0] out233,
  output [WIDTH-1:0] out234,
  output [WIDTH-1:0] out235,
  output [WIDTH-1:0] out236,
  output [WIDTH-1:0] out237,
  output [WIDTH-1:0] out238,
  output [WIDTH-1:0] out239,
  output [WIDTH-1:0] out240,
  output [WIDTH-1:0] out241,
  output [WIDTH-1:0] out242,
  output [WIDTH-1:0] out243,
  output [WIDTH-1:0] out244,
  output [WIDTH-1:0] out245,
  output [WIDTH-1:0] out246,
  output [WIDTH-1:0] out247,
  output [WIDTH-1:0] out248,
  output [WIDTH-1:0] out249,
  output [WIDTH-1:0] out250,
  output [WIDTH-1:0] out251,
  output [WIDTH-1:0] out252,
  output [WIDTH-1:0] out253,
  output [WIDTH-1:0] out254,
  output [WIDTH-1:0] out255
);

  wire [2048-1:0] conf_out;
  wire [WIDTH-1:0] in_reg_wire_0 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_1 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_2 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_3 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_4 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_5 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_6 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_7 [0:256-1];
  wire [64-1:0] net_conf_bus [0:256-1];

  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg0
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus_in),
    .out(net_conf_bus[0])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(1),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_0
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[0]),
    .conf_bus_in(net_conf_bus[0]),
    .swicth_conf_out(conf_out[7:0])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg1
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[0]),
    .out(net_conf_bus[1])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(2),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_1
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[1]),
    .conf_bus_in(net_conf_bus[1]),
    .swicth_conf_out(conf_out[15:8])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[1]),
    .out(net_conf_bus[2])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(3),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_2
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[2]),
    .conf_bus_in(net_conf_bus[2]),
    .swicth_conf_out(conf_out[23:16])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg3
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[2]),
    .out(net_conf_bus[3])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(4),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_3
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[3]),
    .conf_bus_in(net_conf_bus[3]),
    .swicth_conf_out(conf_out[31:24])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg4
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[3]),
    .out(net_conf_bus[4])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(5),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_4
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[4]),
    .conf_bus_in(net_conf_bus[4]),
    .swicth_conf_out(conf_out[39:32])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg5
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[4]),
    .out(net_conf_bus[5])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(6),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_5
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[5]),
    .conf_bus_in(net_conf_bus[5]),
    .swicth_conf_out(conf_out[47:40])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg6
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[5]),
    .out(net_conf_bus[6])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(7),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_6
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[6]),
    .conf_bus_in(net_conf_bus[6]),
    .swicth_conf_out(conf_out[55:48])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg7
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[6]),
    .out(net_conf_bus[7])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(8),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_7
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[7]),
    .conf_bus_in(net_conf_bus[7]),
    .swicth_conf_out(conf_out[63:56])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg8
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[7]),
    .out(net_conf_bus[8])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(9),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_8
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[8]),
    .conf_bus_in(net_conf_bus[8]),
    .swicth_conf_out(conf_out[71:64])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg9
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[8]),
    .out(net_conf_bus[9])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(10),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_9
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[9]),
    .conf_bus_in(net_conf_bus[9]),
    .swicth_conf_out(conf_out[79:72])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg10
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[9]),
    .out(net_conf_bus[10])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(11),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_10
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[10]),
    .conf_bus_in(net_conf_bus[10]),
    .swicth_conf_out(conf_out[87:80])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg11
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[10]),
    .out(net_conf_bus[11])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(12),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_11
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[11]),
    .conf_bus_in(net_conf_bus[11]),
    .swicth_conf_out(conf_out[95:88])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg12
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[11]),
    .out(net_conf_bus[12])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(13),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_12
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[12]),
    .conf_bus_in(net_conf_bus[12]),
    .swicth_conf_out(conf_out[103:96])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg13
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[12]),
    .out(net_conf_bus[13])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(14),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_13
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[13]),
    .conf_bus_in(net_conf_bus[13]),
    .swicth_conf_out(conf_out[111:104])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg14
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[13]),
    .out(net_conf_bus[14])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(15),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_14
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[14]),
    .conf_bus_in(net_conf_bus[14]),
    .swicth_conf_out(conf_out[119:112])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg15
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[14]),
    .out(net_conf_bus[15])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(16),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_15
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[15]),
    .conf_bus_in(net_conf_bus[15]),
    .swicth_conf_out(conf_out[127:120])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg16
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[15]),
    .out(net_conf_bus[16])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(17),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_16
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[16]),
    .conf_bus_in(net_conf_bus[16]),
    .swicth_conf_out(conf_out[135:128])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg17
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[16]),
    .out(net_conf_bus[17])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(18),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_17
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[17]),
    .conf_bus_in(net_conf_bus[17]),
    .swicth_conf_out(conf_out[143:136])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg18
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[17]),
    .out(net_conf_bus[18])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(19),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_18
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[18]),
    .conf_bus_in(net_conf_bus[18]),
    .swicth_conf_out(conf_out[151:144])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg19
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[18]),
    .out(net_conf_bus[19])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(20),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_19
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[19]),
    .conf_bus_in(net_conf_bus[19]),
    .swicth_conf_out(conf_out[159:152])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg20
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[19]),
    .out(net_conf_bus[20])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(21),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_20
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[20]),
    .conf_bus_in(net_conf_bus[20]),
    .swicth_conf_out(conf_out[167:160])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg21
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[20]),
    .out(net_conf_bus[21])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(22),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_21
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[21]),
    .conf_bus_in(net_conf_bus[21]),
    .swicth_conf_out(conf_out[175:168])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg22
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[21]),
    .out(net_conf_bus[22])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(23),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_22
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[22]),
    .conf_bus_in(net_conf_bus[22]),
    .swicth_conf_out(conf_out[183:176])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg23
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[22]),
    .out(net_conf_bus[23])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(24),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_23
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[23]),
    .conf_bus_in(net_conf_bus[23]),
    .swicth_conf_out(conf_out[191:184])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg24
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[23]),
    .out(net_conf_bus[24])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(25),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_24
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[24]),
    .conf_bus_in(net_conf_bus[24]),
    .swicth_conf_out(conf_out[199:192])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg25
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[24]),
    .out(net_conf_bus[25])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(26),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_25
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[25]),
    .conf_bus_in(net_conf_bus[25]),
    .swicth_conf_out(conf_out[207:200])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg26
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[25]),
    .out(net_conf_bus[26])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(27),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_26
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[26]),
    .conf_bus_in(net_conf_bus[26]),
    .swicth_conf_out(conf_out[215:208])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg27
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[26]),
    .out(net_conf_bus[27])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(28),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_27
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[27]),
    .conf_bus_in(net_conf_bus[27]),
    .swicth_conf_out(conf_out[223:216])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg28
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[27]),
    .out(net_conf_bus[28])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(29),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_28
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[28]),
    .conf_bus_in(net_conf_bus[28]),
    .swicth_conf_out(conf_out[231:224])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg29
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[28]),
    .out(net_conf_bus[29])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(30),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_29
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[29]),
    .conf_bus_in(net_conf_bus[29]),
    .swicth_conf_out(conf_out[239:232])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg30
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[29]),
    .out(net_conf_bus[30])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(31),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_30
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[30]),
    .conf_bus_in(net_conf_bus[30]),
    .swicth_conf_out(conf_out[247:240])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg31
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[30]),
    .out(net_conf_bus[31])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(32),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_31
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[31]),
    .conf_bus_in(net_conf_bus[31]),
    .swicth_conf_out(conf_out[255:248])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg32
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[31]),
    .out(net_conf_bus[32])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(33),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_32
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[32]),
    .conf_bus_in(net_conf_bus[32]),
    .swicth_conf_out(conf_out[263:256])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg33
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[32]),
    .out(net_conf_bus[33])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(34),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_33
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[33]),
    .conf_bus_in(net_conf_bus[33]),
    .swicth_conf_out(conf_out[271:264])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg34
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[33]),
    .out(net_conf_bus[34])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(35),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_34
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[34]),
    .conf_bus_in(net_conf_bus[34]),
    .swicth_conf_out(conf_out[279:272])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg35
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[34]),
    .out(net_conf_bus[35])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(36),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_35
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[35]),
    .conf_bus_in(net_conf_bus[35]),
    .swicth_conf_out(conf_out[287:280])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg36
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[35]),
    .out(net_conf_bus[36])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(37),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_36
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[36]),
    .conf_bus_in(net_conf_bus[36]),
    .swicth_conf_out(conf_out[295:288])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg37
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[36]),
    .out(net_conf_bus[37])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(38),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_37
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[37]),
    .conf_bus_in(net_conf_bus[37]),
    .swicth_conf_out(conf_out[303:296])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg38
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[37]),
    .out(net_conf_bus[38])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(39),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_38
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[38]),
    .conf_bus_in(net_conf_bus[38]),
    .swicth_conf_out(conf_out[311:304])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg39
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[38]),
    .out(net_conf_bus[39])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(40),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_39
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[39]),
    .conf_bus_in(net_conf_bus[39]),
    .swicth_conf_out(conf_out[319:312])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg40
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[39]),
    .out(net_conf_bus[40])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(41),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_40
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[40]),
    .conf_bus_in(net_conf_bus[40]),
    .swicth_conf_out(conf_out[327:320])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg41
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[40]),
    .out(net_conf_bus[41])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(42),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_41
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[41]),
    .conf_bus_in(net_conf_bus[41]),
    .swicth_conf_out(conf_out[335:328])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg42
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[41]),
    .out(net_conf_bus[42])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(43),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_42
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[42]),
    .conf_bus_in(net_conf_bus[42]),
    .swicth_conf_out(conf_out[343:336])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg43
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[42]),
    .out(net_conf_bus[43])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(44),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_43
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[43]),
    .conf_bus_in(net_conf_bus[43]),
    .swicth_conf_out(conf_out[351:344])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg44
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[43]),
    .out(net_conf_bus[44])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(45),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_44
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[44]),
    .conf_bus_in(net_conf_bus[44]),
    .swicth_conf_out(conf_out[359:352])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg45
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[44]),
    .out(net_conf_bus[45])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(46),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_45
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[45]),
    .conf_bus_in(net_conf_bus[45]),
    .swicth_conf_out(conf_out[367:360])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg46
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[45]),
    .out(net_conf_bus[46])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(47),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_46
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[46]),
    .conf_bus_in(net_conf_bus[46]),
    .swicth_conf_out(conf_out[375:368])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg47
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[46]),
    .out(net_conf_bus[47])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(48),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_47
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[47]),
    .conf_bus_in(net_conf_bus[47]),
    .swicth_conf_out(conf_out[383:376])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg48
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[47]),
    .out(net_conf_bus[48])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(49),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_48
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[48]),
    .conf_bus_in(net_conf_bus[48]),
    .swicth_conf_out(conf_out[391:384])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg49
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[48]),
    .out(net_conf_bus[49])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(50),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_49
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[49]),
    .conf_bus_in(net_conf_bus[49]),
    .swicth_conf_out(conf_out[399:392])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg50
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[49]),
    .out(net_conf_bus[50])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(51),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_50
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[50]),
    .conf_bus_in(net_conf_bus[50]),
    .swicth_conf_out(conf_out[407:400])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg51
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[50]),
    .out(net_conf_bus[51])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(52),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_51
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[51]),
    .conf_bus_in(net_conf_bus[51]),
    .swicth_conf_out(conf_out[415:408])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg52
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[51]),
    .out(net_conf_bus[52])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(53),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_52
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[52]),
    .conf_bus_in(net_conf_bus[52]),
    .swicth_conf_out(conf_out[423:416])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg53
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[52]),
    .out(net_conf_bus[53])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(54),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_53
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[53]),
    .conf_bus_in(net_conf_bus[53]),
    .swicth_conf_out(conf_out[431:424])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg54
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[53]),
    .out(net_conf_bus[54])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(55),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_54
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[54]),
    .conf_bus_in(net_conf_bus[54]),
    .swicth_conf_out(conf_out[439:432])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg55
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[54]),
    .out(net_conf_bus[55])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(56),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_55
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[55]),
    .conf_bus_in(net_conf_bus[55]),
    .swicth_conf_out(conf_out[447:440])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg56
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[55]),
    .out(net_conf_bus[56])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(57),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_56
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[56]),
    .conf_bus_in(net_conf_bus[56]),
    .swicth_conf_out(conf_out[455:448])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg57
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[56]),
    .out(net_conf_bus[57])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(58),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_57
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[57]),
    .conf_bus_in(net_conf_bus[57]),
    .swicth_conf_out(conf_out[463:456])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg58
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[57]),
    .out(net_conf_bus[58])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(59),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_58
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[58]),
    .conf_bus_in(net_conf_bus[58]),
    .swicth_conf_out(conf_out[471:464])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg59
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[58]),
    .out(net_conf_bus[59])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(60),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_59
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[59]),
    .conf_bus_in(net_conf_bus[59]),
    .swicth_conf_out(conf_out[479:472])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg60
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[59]),
    .out(net_conf_bus[60])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(61),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_60
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[60]),
    .conf_bus_in(net_conf_bus[60]),
    .swicth_conf_out(conf_out[487:480])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg61
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[60]),
    .out(net_conf_bus[61])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(62),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_61
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[61]),
    .conf_bus_in(net_conf_bus[61]),
    .swicth_conf_out(conf_out[495:488])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg62
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[61]),
    .out(net_conf_bus[62])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(63),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_62
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[62]),
    .conf_bus_in(net_conf_bus[62]),
    .swicth_conf_out(conf_out[503:496])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg63
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[62]),
    .out(net_conf_bus[63])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(64),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_63
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[63]),
    .conf_bus_in(net_conf_bus[63]),
    .swicth_conf_out(conf_out[511:504])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg64
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[63]),
    .out(net_conf_bus[64])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(65),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_64
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[64]),
    .conf_bus_in(net_conf_bus[64]),
    .swicth_conf_out(conf_out[519:512])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg65
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[64]),
    .out(net_conf_bus[65])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(66),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_65
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[65]),
    .conf_bus_in(net_conf_bus[65]),
    .swicth_conf_out(conf_out[527:520])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg66
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[65]),
    .out(net_conf_bus[66])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(67),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_66
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[66]),
    .conf_bus_in(net_conf_bus[66]),
    .swicth_conf_out(conf_out[535:528])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg67
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[66]),
    .out(net_conf_bus[67])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(68),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_67
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[67]),
    .conf_bus_in(net_conf_bus[67]),
    .swicth_conf_out(conf_out[543:536])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg68
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[67]),
    .out(net_conf_bus[68])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(69),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_68
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[68]),
    .conf_bus_in(net_conf_bus[68]),
    .swicth_conf_out(conf_out[551:544])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg69
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[68]),
    .out(net_conf_bus[69])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(70),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_69
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[69]),
    .conf_bus_in(net_conf_bus[69]),
    .swicth_conf_out(conf_out[559:552])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg70
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[69]),
    .out(net_conf_bus[70])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(71),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_70
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[70]),
    .conf_bus_in(net_conf_bus[70]),
    .swicth_conf_out(conf_out[567:560])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg71
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[70]),
    .out(net_conf_bus[71])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(72),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_71
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[71]),
    .conf_bus_in(net_conf_bus[71]),
    .swicth_conf_out(conf_out[575:568])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg72
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[71]),
    .out(net_conf_bus[72])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(73),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_72
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[72]),
    .conf_bus_in(net_conf_bus[72]),
    .swicth_conf_out(conf_out[583:576])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg73
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[72]),
    .out(net_conf_bus[73])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(74),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_73
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[73]),
    .conf_bus_in(net_conf_bus[73]),
    .swicth_conf_out(conf_out[591:584])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg74
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[73]),
    .out(net_conf_bus[74])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(75),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_74
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[74]),
    .conf_bus_in(net_conf_bus[74]),
    .swicth_conf_out(conf_out[599:592])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg75
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[74]),
    .out(net_conf_bus[75])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(76),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_75
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[75]),
    .conf_bus_in(net_conf_bus[75]),
    .swicth_conf_out(conf_out[607:600])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg76
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[75]),
    .out(net_conf_bus[76])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(77),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_76
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[76]),
    .conf_bus_in(net_conf_bus[76]),
    .swicth_conf_out(conf_out[615:608])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg77
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[76]),
    .out(net_conf_bus[77])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(78),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_77
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[77]),
    .conf_bus_in(net_conf_bus[77]),
    .swicth_conf_out(conf_out[623:616])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg78
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[77]),
    .out(net_conf_bus[78])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(79),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_78
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[78]),
    .conf_bus_in(net_conf_bus[78]),
    .swicth_conf_out(conf_out[631:624])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg79
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[78]),
    .out(net_conf_bus[79])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(80),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_79
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[79]),
    .conf_bus_in(net_conf_bus[79]),
    .swicth_conf_out(conf_out[639:632])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg80
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[79]),
    .out(net_conf_bus[80])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(81),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_80
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[80]),
    .conf_bus_in(net_conf_bus[80]),
    .swicth_conf_out(conf_out[647:640])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg81
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[80]),
    .out(net_conf_bus[81])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(82),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_81
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[81]),
    .conf_bus_in(net_conf_bus[81]),
    .swicth_conf_out(conf_out[655:648])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg82
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[81]),
    .out(net_conf_bus[82])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(83),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_82
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[82]),
    .conf_bus_in(net_conf_bus[82]),
    .swicth_conf_out(conf_out[663:656])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg83
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[82]),
    .out(net_conf_bus[83])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(84),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_83
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[83]),
    .conf_bus_in(net_conf_bus[83]),
    .swicth_conf_out(conf_out[671:664])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg84
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[83]),
    .out(net_conf_bus[84])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(85),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_84
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[84]),
    .conf_bus_in(net_conf_bus[84]),
    .swicth_conf_out(conf_out[679:672])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg85
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[84]),
    .out(net_conf_bus[85])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(86),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_85
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[85]),
    .conf_bus_in(net_conf_bus[85]),
    .swicth_conf_out(conf_out[687:680])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg86
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[85]),
    .out(net_conf_bus[86])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(87),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_86
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[86]),
    .conf_bus_in(net_conf_bus[86]),
    .swicth_conf_out(conf_out[695:688])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg87
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[86]),
    .out(net_conf_bus[87])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(88),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_87
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[87]),
    .conf_bus_in(net_conf_bus[87]),
    .swicth_conf_out(conf_out[703:696])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg88
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[87]),
    .out(net_conf_bus[88])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(89),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_88
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[88]),
    .conf_bus_in(net_conf_bus[88]),
    .swicth_conf_out(conf_out[711:704])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg89
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[88]),
    .out(net_conf_bus[89])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(90),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_89
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[89]),
    .conf_bus_in(net_conf_bus[89]),
    .swicth_conf_out(conf_out[719:712])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg90
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[89]),
    .out(net_conf_bus[90])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(91),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_90
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[90]),
    .conf_bus_in(net_conf_bus[90]),
    .swicth_conf_out(conf_out[727:720])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg91
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[90]),
    .out(net_conf_bus[91])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(92),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_91
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[91]),
    .conf_bus_in(net_conf_bus[91]),
    .swicth_conf_out(conf_out[735:728])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg92
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[91]),
    .out(net_conf_bus[92])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(93),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_92
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[92]),
    .conf_bus_in(net_conf_bus[92]),
    .swicth_conf_out(conf_out[743:736])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg93
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[92]),
    .out(net_conf_bus[93])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(94),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_93
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[93]),
    .conf_bus_in(net_conf_bus[93]),
    .swicth_conf_out(conf_out[751:744])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg94
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[93]),
    .out(net_conf_bus[94])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(95),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_94
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[94]),
    .conf_bus_in(net_conf_bus[94]),
    .swicth_conf_out(conf_out[759:752])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg95
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[94]),
    .out(net_conf_bus[95])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(96),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_95
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[95]),
    .conf_bus_in(net_conf_bus[95]),
    .swicth_conf_out(conf_out[767:760])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg96
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[95]),
    .out(net_conf_bus[96])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(97),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_96
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[96]),
    .conf_bus_in(net_conf_bus[96]),
    .swicth_conf_out(conf_out[775:768])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg97
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[96]),
    .out(net_conf_bus[97])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(98),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_97
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[97]),
    .conf_bus_in(net_conf_bus[97]),
    .swicth_conf_out(conf_out[783:776])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg98
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[97]),
    .out(net_conf_bus[98])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(99),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_98
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[98]),
    .conf_bus_in(net_conf_bus[98]),
    .swicth_conf_out(conf_out[791:784])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg99
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[98]),
    .out(net_conf_bus[99])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(100),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_99
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[99]),
    .conf_bus_in(net_conf_bus[99]),
    .swicth_conf_out(conf_out[799:792])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg100
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[99]),
    .out(net_conf_bus[100])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(101),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_100
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[100]),
    .conf_bus_in(net_conf_bus[100]),
    .swicth_conf_out(conf_out[807:800])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg101
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[100]),
    .out(net_conf_bus[101])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(102),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_101
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[101]),
    .conf_bus_in(net_conf_bus[101]),
    .swicth_conf_out(conf_out[815:808])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg102
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[101]),
    .out(net_conf_bus[102])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(103),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_102
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[102]),
    .conf_bus_in(net_conf_bus[102]),
    .swicth_conf_out(conf_out[823:816])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg103
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[102]),
    .out(net_conf_bus[103])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(104),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_103
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[103]),
    .conf_bus_in(net_conf_bus[103]),
    .swicth_conf_out(conf_out[831:824])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg104
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[103]),
    .out(net_conf_bus[104])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(105),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_104
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[104]),
    .conf_bus_in(net_conf_bus[104]),
    .swicth_conf_out(conf_out[839:832])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg105
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[104]),
    .out(net_conf_bus[105])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(106),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_105
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[105]),
    .conf_bus_in(net_conf_bus[105]),
    .swicth_conf_out(conf_out[847:840])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg106
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[105]),
    .out(net_conf_bus[106])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(107),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_106
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[106]),
    .conf_bus_in(net_conf_bus[106]),
    .swicth_conf_out(conf_out[855:848])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg107
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[106]),
    .out(net_conf_bus[107])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(108),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_107
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[107]),
    .conf_bus_in(net_conf_bus[107]),
    .swicth_conf_out(conf_out[863:856])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg108
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[107]),
    .out(net_conf_bus[108])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(109),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_108
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[108]),
    .conf_bus_in(net_conf_bus[108]),
    .swicth_conf_out(conf_out[871:864])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg109
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[108]),
    .out(net_conf_bus[109])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(110),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_109
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[109]),
    .conf_bus_in(net_conf_bus[109]),
    .swicth_conf_out(conf_out[879:872])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg110
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[109]),
    .out(net_conf_bus[110])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(111),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_110
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[110]),
    .conf_bus_in(net_conf_bus[110]),
    .swicth_conf_out(conf_out[887:880])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg111
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[110]),
    .out(net_conf_bus[111])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(112),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_111
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[111]),
    .conf_bus_in(net_conf_bus[111]),
    .swicth_conf_out(conf_out[895:888])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg112
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[111]),
    .out(net_conf_bus[112])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(113),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_112
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[112]),
    .conf_bus_in(net_conf_bus[112]),
    .swicth_conf_out(conf_out[903:896])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg113
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[112]),
    .out(net_conf_bus[113])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(114),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_113
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[113]),
    .conf_bus_in(net_conf_bus[113]),
    .swicth_conf_out(conf_out[911:904])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg114
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[113]),
    .out(net_conf_bus[114])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(115),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_114
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[114]),
    .conf_bus_in(net_conf_bus[114]),
    .swicth_conf_out(conf_out[919:912])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg115
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[114]),
    .out(net_conf_bus[115])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(116),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_115
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[115]),
    .conf_bus_in(net_conf_bus[115]),
    .swicth_conf_out(conf_out[927:920])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg116
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[115]),
    .out(net_conf_bus[116])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(117),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_116
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[116]),
    .conf_bus_in(net_conf_bus[116]),
    .swicth_conf_out(conf_out[935:928])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg117
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[116]),
    .out(net_conf_bus[117])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(118),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_117
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[117]),
    .conf_bus_in(net_conf_bus[117]),
    .swicth_conf_out(conf_out[943:936])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg118
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[117]),
    .out(net_conf_bus[118])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(119),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_118
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[118]),
    .conf_bus_in(net_conf_bus[118]),
    .swicth_conf_out(conf_out[951:944])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg119
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[118]),
    .out(net_conf_bus[119])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(120),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_119
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[119]),
    .conf_bus_in(net_conf_bus[119]),
    .swicth_conf_out(conf_out[959:952])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg120
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[119]),
    .out(net_conf_bus[120])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(121),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_120
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[120]),
    .conf_bus_in(net_conf_bus[120]),
    .swicth_conf_out(conf_out[967:960])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg121
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[120]),
    .out(net_conf_bus[121])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(122),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_121
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[121]),
    .conf_bus_in(net_conf_bus[121]),
    .swicth_conf_out(conf_out[975:968])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg122
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[121]),
    .out(net_conf_bus[122])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(123),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_122
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[122]),
    .conf_bus_in(net_conf_bus[122]),
    .swicth_conf_out(conf_out[983:976])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg123
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[122]),
    .out(net_conf_bus[123])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(124),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_123
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[123]),
    .conf_bus_in(net_conf_bus[123]),
    .swicth_conf_out(conf_out[991:984])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg124
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[123]),
    .out(net_conf_bus[124])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(125),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_124
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[124]),
    .conf_bus_in(net_conf_bus[124]),
    .swicth_conf_out(conf_out[999:992])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg125
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[124]),
    .out(net_conf_bus[125])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(126),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_125
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[125]),
    .conf_bus_in(net_conf_bus[125]),
    .swicth_conf_out(conf_out[1007:1000])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg126
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[125]),
    .out(net_conf_bus[126])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(127),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_126
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[126]),
    .conf_bus_in(net_conf_bus[126]),
    .swicth_conf_out(conf_out[1015:1008])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg127
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[126]),
    .out(net_conf_bus[127])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(128),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_127
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[127]),
    .conf_bus_in(net_conf_bus[127]),
    .swicth_conf_out(conf_out[1023:1016])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg128
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[127]),
    .out(net_conf_bus[128])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(129),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_128
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[128]),
    .conf_bus_in(net_conf_bus[128]),
    .swicth_conf_out(conf_out[1031:1024])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg129
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[128]),
    .out(net_conf_bus[129])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(130),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_129
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[129]),
    .conf_bus_in(net_conf_bus[129]),
    .swicth_conf_out(conf_out[1039:1032])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg130
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[129]),
    .out(net_conf_bus[130])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(131),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_130
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[130]),
    .conf_bus_in(net_conf_bus[130]),
    .swicth_conf_out(conf_out[1047:1040])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg131
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[130]),
    .out(net_conf_bus[131])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(132),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_131
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[131]),
    .conf_bus_in(net_conf_bus[131]),
    .swicth_conf_out(conf_out[1055:1048])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg132
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[131]),
    .out(net_conf_bus[132])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(133),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_132
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[132]),
    .conf_bus_in(net_conf_bus[132]),
    .swicth_conf_out(conf_out[1063:1056])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg133
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[132]),
    .out(net_conf_bus[133])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(134),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_133
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[133]),
    .conf_bus_in(net_conf_bus[133]),
    .swicth_conf_out(conf_out[1071:1064])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg134
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[133]),
    .out(net_conf_bus[134])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(135),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_134
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[134]),
    .conf_bus_in(net_conf_bus[134]),
    .swicth_conf_out(conf_out[1079:1072])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg135
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[134]),
    .out(net_conf_bus[135])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(136),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_135
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[135]),
    .conf_bus_in(net_conf_bus[135]),
    .swicth_conf_out(conf_out[1087:1080])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg136
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[135]),
    .out(net_conf_bus[136])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(137),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_136
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[136]),
    .conf_bus_in(net_conf_bus[136]),
    .swicth_conf_out(conf_out[1095:1088])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg137
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[136]),
    .out(net_conf_bus[137])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(138),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_137
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[137]),
    .conf_bus_in(net_conf_bus[137]),
    .swicth_conf_out(conf_out[1103:1096])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg138
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[137]),
    .out(net_conf_bus[138])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(139),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_138
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[138]),
    .conf_bus_in(net_conf_bus[138]),
    .swicth_conf_out(conf_out[1111:1104])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg139
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[138]),
    .out(net_conf_bus[139])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(140),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_139
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[139]),
    .conf_bus_in(net_conf_bus[139]),
    .swicth_conf_out(conf_out[1119:1112])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg140
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[139]),
    .out(net_conf_bus[140])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(141),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_140
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[140]),
    .conf_bus_in(net_conf_bus[140]),
    .swicth_conf_out(conf_out[1127:1120])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg141
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[140]),
    .out(net_conf_bus[141])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(142),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_141
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[141]),
    .conf_bus_in(net_conf_bus[141]),
    .swicth_conf_out(conf_out[1135:1128])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg142
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[141]),
    .out(net_conf_bus[142])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(143),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_142
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[142]),
    .conf_bus_in(net_conf_bus[142]),
    .swicth_conf_out(conf_out[1143:1136])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg143
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[142]),
    .out(net_conf_bus[143])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(144),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_143
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[143]),
    .conf_bus_in(net_conf_bus[143]),
    .swicth_conf_out(conf_out[1151:1144])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg144
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[143]),
    .out(net_conf_bus[144])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(145),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_144
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[144]),
    .conf_bus_in(net_conf_bus[144]),
    .swicth_conf_out(conf_out[1159:1152])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg145
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[144]),
    .out(net_conf_bus[145])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(146),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_145
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[145]),
    .conf_bus_in(net_conf_bus[145]),
    .swicth_conf_out(conf_out[1167:1160])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg146
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[145]),
    .out(net_conf_bus[146])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(147),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_146
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[146]),
    .conf_bus_in(net_conf_bus[146]),
    .swicth_conf_out(conf_out[1175:1168])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg147
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[146]),
    .out(net_conf_bus[147])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(148),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_147
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[147]),
    .conf_bus_in(net_conf_bus[147]),
    .swicth_conf_out(conf_out[1183:1176])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg148
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[147]),
    .out(net_conf_bus[148])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(149),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_148
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[148]),
    .conf_bus_in(net_conf_bus[148]),
    .swicth_conf_out(conf_out[1191:1184])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg149
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[148]),
    .out(net_conf_bus[149])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(150),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_149
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[149]),
    .conf_bus_in(net_conf_bus[149]),
    .swicth_conf_out(conf_out[1199:1192])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg150
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[149]),
    .out(net_conf_bus[150])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(151),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_150
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[150]),
    .conf_bus_in(net_conf_bus[150]),
    .swicth_conf_out(conf_out[1207:1200])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg151
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[150]),
    .out(net_conf_bus[151])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(152),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_151
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[151]),
    .conf_bus_in(net_conf_bus[151]),
    .swicth_conf_out(conf_out[1215:1208])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg152
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[151]),
    .out(net_conf_bus[152])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(153),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_152
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[152]),
    .conf_bus_in(net_conf_bus[152]),
    .swicth_conf_out(conf_out[1223:1216])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg153
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[152]),
    .out(net_conf_bus[153])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(154),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_153
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[153]),
    .conf_bus_in(net_conf_bus[153]),
    .swicth_conf_out(conf_out[1231:1224])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg154
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[153]),
    .out(net_conf_bus[154])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(155),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_154
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[154]),
    .conf_bus_in(net_conf_bus[154]),
    .swicth_conf_out(conf_out[1239:1232])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg155
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[154]),
    .out(net_conf_bus[155])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(156),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_155
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[155]),
    .conf_bus_in(net_conf_bus[155]),
    .swicth_conf_out(conf_out[1247:1240])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg156
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[155]),
    .out(net_conf_bus[156])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(157),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_156
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[156]),
    .conf_bus_in(net_conf_bus[156]),
    .swicth_conf_out(conf_out[1255:1248])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg157
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[156]),
    .out(net_conf_bus[157])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(158),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_157
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[157]),
    .conf_bus_in(net_conf_bus[157]),
    .swicth_conf_out(conf_out[1263:1256])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg158
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[157]),
    .out(net_conf_bus[158])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(159),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_158
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[158]),
    .conf_bus_in(net_conf_bus[158]),
    .swicth_conf_out(conf_out[1271:1264])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg159
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[158]),
    .out(net_conf_bus[159])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(160),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_159
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[159]),
    .conf_bus_in(net_conf_bus[159]),
    .swicth_conf_out(conf_out[1279:1272])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg160
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[159]),
    .out(net_conf_bus[160])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(161),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_160
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[160]),
    .conf_bus_in(net_conf_bus[160]),
    .swicth_conf_out(conf_out[1287:1280])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg161
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[160]),
    .out(net_conf_bus[161])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(162),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_161
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[161]),
    .conf_bus_in(net_conf_bus[161]),
    .swicth_conf_out(conf_out[1295:1288])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg162
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[161]),
    .out(net_conf_bus[162])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(163),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_162
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[162]),
    .conf_bus_in(net_conf_bus[162]),
    .swicth_conf_out(conf_out[1303:1296])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg163
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[162]),
    .out(net_conf_bus[163])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(164),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_163
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[163]),
    .conf_bus_in(net_conf_bus[163]),
    .swicth_conf_out(conf_out[1311:1304])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg164
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[163]),
    .out(net_conf_bus[164])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(165),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_164
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[164]),
    .conf_bus_in(net_conf_bus[164]),
    .swicth_conf_out(conf_out[1319:1312])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg165
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[164]),
    .out(net_conf_bus[165])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(166),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_165
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[165]),
    .conf_bus_in(net_conf_bus[165]),
    .swicth_conf_out(conf_out[1327:1320])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg166
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[165]),
    .out(net_conf_bus[166])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(167),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_166
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[166]),
    .conf_bus_in(net_conf_bus[166]),
    .swicth_conf_out(conf_out[1335:1328])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg167
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[166]),
    .out(net_conf_bus[167])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(168),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_167
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[167]),
    .conf_bus_in(net_conf_bus[167]),
    .swicth_conf_out(conf_out[1343:1336])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg168
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[167]),
    .out(net_conf_bus[168])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(169),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_168
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[168]),
    .conf_bus_in(net_conf_bus[168]),
    .swicth_conf_out(conf_out[1351:1344])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg169
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[168]),
    .out(net_conf_bus[169])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(170),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_169
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[169]),
    .conf_bus_in(net_conf_bus[169]),
    .swicth_conf_out(conf_out[1359:1352])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg170
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[169]),
    .out(net_conf_bus[170])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(171),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_170
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[170]),
    .conf_bus_in(net_conf_bus[170]),
    .swicth_conf_out(conf_out[1367:1360])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg171
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[170]),
    .out(net_conf_bus[171])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(172),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_171
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[171]),
    .conf_bus_in(net_conf_bus[171]),
    .swicth_conf_out(conf_out[1375:1368])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg172
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[171]),
    .out(net_conf_bus[172])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(173),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_172
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[172]),
    .conf_bus_in(net_conf_bus[172]),
    .swicth_conf_out(conf_out[1383:1376])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg173
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[172]),
    .out(net_conf_bus[173])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(174),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_173
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[173]),
    .conf_bus_in(net_conf_bus[173]),
    .swicth_conf_out(conf_out[1391:1384])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg174
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[173]),
    .out(net_conf_bus[174])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(175),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_174
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[174]),
    .conf_bus_in(net_conf_bus[174]),
    .swicth_conf_out(conf_out[1399:1392])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg175
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[174]),
    .out(net_conf_bus[175])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(176),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_175
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[175]),
    .conf_bus_in(net_conf_bus[175]),
    .swicth_conf_out(conf_out[1407:1400])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg176
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[175]),
    .out(net_conf_bus[176])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(177),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_176
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[176]),
    .conf_bus_in(net_conf_bus[176]),
    .swicth_conf_out(conf_out[1415:1408])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg177
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[176]),
    .out(net_conf_bus[177])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(178),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_177
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[177]),
    .conf_bus_in(net_conf_bus[177]),
    .swicth_conf_out(conf_out[1423:1416])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg178
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[177]),
    .out(net_conf_bus[178])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(179),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_178
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[178]),
    .conf_bus_in(net_conf_bus[178]),
    .swicth_conf_out(conf_out[1431:1424])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg179
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[178]),
    .out(net_conf_bus[179])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(180),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_179
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[179]),
    .conf_bus_in(net_conf_bus[179]),
    .swicth_conf_out(conf_out[1439:1432])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg180
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[179]),
    .out(net_conf_bus[180])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(181),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_180
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[180]),
    .conf_bus_in(net_conf_bus[180]),
    .swicth_conf_out(conf_out[1447:1440])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg181
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[180]),
    .out(net_conf_bus[181])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(182),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_181
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[181]),
    .conf_bus_in(net_conf_bus[181]),
    .swicth_conf_out(conf_out[1455:1448])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg182
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[181]),
    .out(net_conf_bus[182])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(183),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_182
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[182]),
    .conf_bus_in(net_conf_bus[182]),
    .swicth_conf_out(conf_out[1463:1456])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg183
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[182]),
    .out(net_conf_bus[183])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(184),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_183
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[183]),
    .conf_bus_in(net_conf_bus[183]),
    .swicth_conf_out(conf_out[1471:1464])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg184
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[183]),
    .out(net_conf_bus[184])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(185),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_184
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[184]),
    .conf_bus_in(net_conf_bus[184]),
    .swicth_conf_out(conf_out[1479:1472])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg185
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[184]),
    .out(net_conf_bus[185])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(186),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_185
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[185]),
    .conf_bus_in(net_conf_bus[185]),
    .swicth_conf_out(conf_out[1487:1480])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg186
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[185]),
    .out(net_conf_bus[186])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(187),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_186
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[186]),
    .conf_bus_in(net_conf_bus[186]),
    .swicth_conf_out(conf_out[1495:1488])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg187
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[186]),
    .out(net_conf_bus[187])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(188),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_187
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[187]),
    .conf_bus_in(net_conf_bus[187]),
    .swicth_conf_out(conf_out[1503:1496])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg188
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[187]),
    .out(net_conf_bus[188])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(189),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_188
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[188]),
    .conf_bus_in(net_conf_bus[188]),
    .swicth_conf_out(conf_out[1511:1504])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg189
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[188]),
    .out(net_conf_bus[189])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(190),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_189
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[189]),
    .conf_bus_in(net_conf_bus[189]),
    .swicth_conf_out(conf_out[1519:1512])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg190
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[189]),
    .out(net_conf_bus[190])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(191),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_190
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[190]),
    .conf_bus_in(net_conf_bus[190]),
    .swicth_conf_out(conf_out[1527:1520])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg191
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[190]),
    .out(net_conf_bus[191])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(192),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_191
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[191]),
    .conf_bus_in(net_conf_bus[191]),
    .swicth_conf_out(conf_out[1535:1528])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg192
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[191]),
    .out(net_conf_bus[192])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(193),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_192
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[192]),
    .conf_bus_in(net_conf_bus[192]),
    .swicth_conf_out(conf_out[1543:1536])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg193
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[192]),
    .out(net_conf_bus[193])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(194),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_193
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[193]),
    .conf_bus_in(net_conf_bus[193]),
    .swicth_conf_out(conf_out[1551:1544])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg194
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[193]),
    .out(net_conf_bus[194])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(195),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_194
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[194]),
    .conf_bus_in(net_conf_bus[194]),
    .swicth_conf_out(conf_out[1559:1552])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg195
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[194]),
    .out(net_conf_bus[195])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(196),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_195
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[195]),
    .conf_bus_in(net_conf_bus[195]),
    .swicth_conf_out(conf_out[1567:1560])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg196
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[195]),
    .out(net_conf_bus[196])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(197),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_196
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[196]),
    .conf_bus_in(net_conf_bus[196]),
    .swicth_conf_out(conf_out[1575:1568])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg197
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[196]),
    .out(net_conf_bus[197])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(198),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_197
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[197]),
    .conf_bus_in(net_conf_bus[197]),
    .swicth_conf_out(conf_out[1583:1576])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg198
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[197]),
    .out(net_conf_bus[198])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(199),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_198
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[198]),
    .conf_bus_in(net_conf_bus[198]),
    .swicth_conf_out(conf_out[1591:1584])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg199
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[198]),
    .out(net_conf_bus[199])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(200),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_199
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[199]),
    .conf_bus_in(net_conf_bus[199]),
    .swicth_conf_out(conf_out[1599:1592])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg200
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[199]),
    .out(net_conf_bus[200])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(201),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_200
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[200]),
    .conf_bus_in(net_conf_bus[200]),
    .swicth_conf_out(conf_out[1607:1600])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg201
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[200]),
    .out(net_conf_bus[201])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(202),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_201
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[201]),
    .conf_bus_in(net_conf_bus[201]),
    .swicth_conf_out(conf_out[1615:1608])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg202
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[201]),
    .out(net_conf_bus[202])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(203),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_202
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[202]),
    .conf_bus_in(net_conf_bus[202]),
    .swicth_conf_out(conf_out[1623:1616])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg203
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[202]),
    .out(net_conf_bus[203])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(204),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_203
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[203]),
    .conf_bus_in(net_conf_bus[203]),
    .swicth_conf_out(conf_out[1631:1624])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg204
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[203]),
    .out(net_conf_bus[204])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(205),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_204
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[204]),
    .conf_bus_in(net_conf_bus[204]),
    .swicth_conf_out(conf_out[1639:1632])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg205
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[204]),
    .out(net_conf_bus[205])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(206),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_205
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[205]),
    .conf_bus_in(net_conf_bus[205]),
    .swicth_conf_out(conf_out[1647:1640])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg206
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[205]),
    .out(net_conf_bus[206])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(207),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_206
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[206]),
    .conf_bus_in(net_conf_bus[206]),
    .swicth_conf_out(conf_out[1655:1648])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg207
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[206]),
    .out(net_conf_bus[207])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(208),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_207
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[207]),
    .conf_bus_in(net_conf_bus[207]),
    .swicth_conf_out(conf_out[1663:1656])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg208
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[207]),
    .out(net_conf_bus[208])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(209),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_208
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[208]),
    .conf_bus_in(net_conf_bus[208]),
    .swicth_conf_out(conf_out[1671:1664])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg209
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[208]),
    .out(net_conf_bus[209])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(210),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_209
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[209]),
    .conf_bus_in(net_conf_bus[209]),
    .swicth_conf_out(conf_out[1679:1672])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg210
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[209]),
    .out(net_conf_bus[210])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(211),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_210
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[210]),
    .conf_bus_in(net_conf_bus[210]),
    .swicth_conf_out(conf_out[1687:1680])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg211
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[210]),
    .out(net_conf_bus[211])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(212),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_211
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[211]),
    .conf_bus_in(net_conf_bus[211]),
    .swicth_conf_out(conf_out[1695:1688])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg212
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[211]),
    .out(net_conf_bus[212])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(213),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_212
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[212]),
    .conf_bus_in(net_conf_bus[212]),
    .swicth_conf_out(conf_out[1703:1696])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg213
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[212]),
    .out(net_conf_bus[213])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(214),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_213
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[213]),
    .conf_bus_in(net_conf_bus[213]),
    .swicth_conf_out(conf_out[1711:1704])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg214
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[213]),
    .out(net_conf_bus[214])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(215),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_214
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[214]),
    .conf_bus_in(net_conf_bus[214]),
    .swicth_conf_out(conf_out[1719:1712])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg215
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[214]),
    .out(net_conf_bus[215])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(216),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_215
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[215]),
    .conf_bus_in(net_conf_bus[215]),
    .swicth_conf_out(conf_out[1727:1720])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg216
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[215]),
    .out(net_conf_bus[216])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(217),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_216
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[216]),
    .conf_bus_in(net_conf_bus[216]),
    .swicth_conf_out(conf_out[1735:1728])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg217
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[216]),
    .out(net_conf_bus[217])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(218),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_217
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[217]),
    .conf_bus_in(net_conf_bus[217]),
    .swicth_conf_out(conf_out[1743:1736])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg218
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[217]),
    .out(net_conf_bus[218])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(219),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_218
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[218]),
    .conf_bus_in(net_conf_bus[218]),
    .swicth_conf_out(conf_out[1751:1744])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg219
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[218]),
    .out(net_conf_bus[219])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(220),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_219
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[219]),
    .conf_bus_in(net_conf_bus[219]),
    .swicth_conf_out(conf_out[1759:1752])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg220
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[219]),
    .out(net_conf_bus[220])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(221),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_220
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[220]),
    .conf_bus_in(net_conf_bus[220]),
    .swicth_conf_out(conf_out[1767:1760])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg221
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[220]),
    .out(net_conf_bus[221])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(222),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_221
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[221]),
    .conf_bus_in(net_conf_bus[221]),
    .swicth_conf_out(conf_out[1775:1768])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg222
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[221]),
    .out(net_conf_bus[222])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(223),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_222
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[222]),
    .conf_bus_in(net_conf_bus[222]),
    .swicth_conf_out(conf_out[1783:1776])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg223
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[222]),
    .out(net_conf_bus[223])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(224),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_223
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[223]),
    .conf_bus_in(net_conf_bus[223]),
    .swicth_conf_out(conf_out[1791:1784])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg224
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[223]),
    .out(net_conf_bus[224])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(225),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_224
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[224]),
    .conf_bus_in(net_conf_bus[224]),
    .swicth_conf_out(conf_out[1799:1792])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg225
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[224]),
    .out(net_conf_bus[225])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(226),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_225
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[225]),
    .conf_bus_in(net_conf_bus[225]),
    .swicth_conf_out(conf_out[1807:1800])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg226
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[225]),
    .out(net_conf_bus[226])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(227),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_226
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[226]),
    .conf_bus_in(net_conf_bus[226]),
    .swicth_conf_out(conf_out[1815:1808])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg227
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[226]),
    .out(net_conf_bus[227])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(228),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_227
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[227]),
    .conf_bus_in(net_conf_bus[227]),
    .swicth_conf_out(conf_out[1823:1816])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg228
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[227]),
    .out(net_conf_bus[228])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(229),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_228
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[228]),
    .conf_bus_in(net_conf_bus[228]),
    .swicth_conf_out(conf_out[1831:1824])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg229
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[228]),
    .out(net_conf_bus[229])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(230),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_229
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[229]),
    .conf_bus_in(net_conf_bus[229]),
    .swicth_conf_out(conf_out[1839:1832])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg230
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[229]),
    .out(net_conf_bus[230])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(231),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_230
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[230]),
    .conf_bus_in(net_conf_bus[230]),
    .swicth_conf_out(conf_out[1847:1840])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg231
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[230]),
    .out(net_conf_bus[231])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(232),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_231
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[231]),
    .conf_bus_in(net_conf_bus[231]),
    .swicth_conf_out(conf_out[1855:1848])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg232
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[231]),
    .out(net_conf_bus[232])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(233),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_232
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[232]),
    .conf_bus_in(net_conf_bus[232]),
    .swicth_conf_out(conf_out[1863:1856])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg233
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[232]),
    .out(net_conf_bus[233])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(234),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_233
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[233]),
    .conf_bus_in(net_conf_bus[233]),
    .swicth_conf_out(conf_out[1871:1864])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg234
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[233]),
    .out(net_conf_bus[234])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(235),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_234
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[234]),
    .conf_bus_in(net_conf_bus[234]),
    .swicth_conf_out(conf_out[1879:1872])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg235
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[234]),
    .out(net_conf_bus[235])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(236),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_235
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[235]),
    .conf_bus_in(net_conf_bus[235]),
    .swicth_conf_out(conf_out[1887:1880])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg236
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[235]),
    .out(net_conf_bus[236])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(237),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_236
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[236]),
    .conf_bus_in(net_conf_bus[236]),
    .swicth_conf_out(conf_out[1895:1888])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg237
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[236]),
    .out(net_conf_bus[237])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(238),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_237
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[237]),
    .conf_bus_in(net_conf_bus[237]),
    .swicth_conf_out(conf_out[1903:1896])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg238
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[237]),
    .out(net_conf_bus[238])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(239),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_238
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[238]),
    .conf_bus_in(net_conf_bus[238]),
    .swicth_conf_out(conf_out[1911:1904])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg239
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[238]),
    .out(net_conf_bus[239])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(240),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_239
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[239]),
    .conf_bus_in(net_conf_bus[239]),
    .swicth_conf_out(conf_out[1919:1912])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg240
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[239]),
    .out(net_conf_bus[240])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(241),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_240
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[240]),
    .conf_bus_in(net_conf_bus[240]),
    .swicth_conf_out(conf_out[1927:1920])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg241
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[240]),
    .out(net_conf_bus[241])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(242),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_241
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[241]),
    .conf_bus_in(net_conf_bus[241]),
    .swicth_conf_out(conf_out[1935:1928])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg242
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[241]),
    .out(net_conf_bus[242])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(243),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_242
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[242]),
    .conf_bus_in(net_conf_bus[242]),
    .swicth_conf_out(conf_out[1943:1936])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg243
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[242]),
    .out(net_conf_bus[243])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(244),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_243
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[243]),
    .conf_bus_in(net_conf_bus[243]),
    .swicth_conf_out(conf_out[1951:1944])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg244
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[243]),
    .out(net_conf_bus[244])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(245),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_244
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[244]),
    .conf_bus_in(net_conf_bus[244]),
    .swicth_conf_out(conf_out[1959:1952])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg245
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[244]),
    .out(net_conf_bus[245])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(246),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_245
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[245]),
    .conf_bus_in(net_conf_bus[245]),
    .swicth_conf_out(conf_out[1967:1960])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg246
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[245]),
    .out(net_conf_bus[246])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(247),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_246
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[246]),
    .conf_bus_in(net_conf_bus[246]),
    .swicth_conf_out(conf_out[1975:1968])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg247
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[246]),
    .out(net_conf_bus[247])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(248),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_247
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[247]),
    .conf_bus_in(net_conf_bus[247]),
    .swicth_conf_out(conf_out[1983:1976])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg248
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[247]),
    .out(net_conf_bus[248])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(249),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_248
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[248]),
    .conf_bus_in(net_conf_bus[248]),
    .swicth_conf_out(conf_out[1991:1984])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg249
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[248]),
    .out(net_conf_bus[249])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(250),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_249
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[249]),
    .conf_bus_in(net_conf_bus[249]),
    .swicth_conf_out(conf_out[1999:1992])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg250
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[249]),
    .out(net_conf_bus[250])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(251),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_250
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[250]),
    .conf_bus_in(net_conf_bus[250]),
    .swicth_conf_out(conf_out[2007:2000])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg251
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[250]),
    .out(net_conf_bus[251])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(252),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_251
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[251]),
    .conf_bus_in(net_conf_bus[251]),
    .swicth_conf_out(conf_out[2015:2008])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg252
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[251]),
    .out(net_conf_bus[252])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(253),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_252
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[252]),
    .conf_bus_in(net_conf_bus[252]),
    .swicth_conf_out(conf_out[2023:2016])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg253
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[252]),
    .out(net_conf_bus[253])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(254),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_253
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[253]),
    .conf_bus_in(net_conf_bus[253]),
    .swicth_conf_out(conf_out[2031:2024])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg254
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[253]),
    .out(net_conf_bus[254])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(255),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_254
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[254]),
    .conf_bus_in(net_conf_bus[254]),
    .swicth_conf_out(conf_out[2039:2032])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg255
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[254]),
    .out(net_conf_bus[255])
  );


  swicth_conf_control_8_8
  #(
    .SWICTH_NUMBER(256),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_255
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en_pc_net[255]),
    .conf_bus_in(net_conf_bus[255]),
    .swicth_conf_out(conf_out[2047:2040])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[0]),
    .in(in0),
    .out(in_reg_wire_0[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1]),
    .in(in1),
    .out(in_reg_wire_0[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[2]),
    .in(in2),
    .out(in_reg_wire_0[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[3]),
    .in(in3),
    .out(in_reg_wire_0[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[4]),
    .in(in4),
    .out(in_reg_wire_0[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[5]),
    .in(in5),
    .out(in_reg_wire_0[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[6]),
    .in(in6),
    .out(in_reg_wire_0[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[7]),
    .in(in7),
    .out(in_reg_wire_0[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[8]),
    .in(in8),
    .out(in_reg_wire_0[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[9]),
    .in(in9),
    .out(in_reg_wire_0[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[10]),
    .in(in10),
    .out(in_reg_wire_0[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[11]),
    .in(in11),
    .out(in_reg_wire_0[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[12]),
    .in(in12),
    .out(in_reg_wire_0[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[13]),
    .in(in13),
    .out(in_reg_wire_0[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[14]),
    .in(in14),
    .out(in_reg_wire_0[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[15]),
    .in(in15),
    .out(in_reg_wire_0[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[16]),
    .in(in16),
    .out(in_reg_wire_0[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[17]),
    .in(in17),
    .out(in_reg_wire_0[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[18]),
    .in(in18),
    .out(in_reg_wire_0[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[19]),
    .in(in19),
    .out(in_reg_wire_0[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[20]),
    .in(in20),
    .out(in_reg_wire_0[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[21]),
    .in(in21),
    .out(in_reg_wire_0[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[22]),
    .in(in22),
    .out(in_reg_wire_0[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[23]),
    .in(in23),
    .out(in_reg_wire_0[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[24]),
    .in(in24),
    .out(in_reg_wire_0[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[25]),
    .in(in25),
    .out(in_reg_wire_0[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[26]),
    .in(in26),
    .out(in_reg_wire_0[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[27]),
    .in(in27),
    .out(in_reg_wire_0[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[28]),
    .in(in28),
    .out(in_reg_wire_0[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[29]),
    .in(in29),
    .out(in_reg_wire_0[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[30]),
    .in(in30),
    .out(in_reg_wire_0[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[31]),
    .in(in31),
    .out(in_reg_wire_0[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[32]),
    .in(in32),
    .out(in_reg_wire_0[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[33]),
    .in(in33),
    .out(in_reg_wire_0[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[34]),
    .in(in34),
    .out(in_reg_wire_0[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[35]),
    .in(in35),
    .out(in_reg_wire_0[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[36]),
    .in(in36),
    .out(in_reg_wire_0[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[37]),
    .in(in37),
    .out(in_reg_wire_0[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[38]),
    .in(in38),
    .out(in_reg_wire_0[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[39]),
    .in(in39),
    .out(in_reg_wire_0[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[40]),
    .in(in40),
    .out(in_reg_wire_0[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[41]),
    .in(in41),
    .out(in_reg_wire_0[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[42]),
    .in(in42),
    .out(in_reg_wire_0[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[43]),
    .in(in43),
    .out(in_reg_wire_0[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[44]),
    .in(in44),
    .out(in_reg_wire_0[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[45]),
    .in(in45),
    .out(in_reg_wire_0[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[46]),
    .in(in46),
    .out(in_reg_wire_0[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[47]),
    .in(in47),
    .out(in_reg_wire_0[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[48]),
    .in(in48),
    .out(in_reg_wire_0[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[49]),
    .in(in49),
    .out(in_reg_wire_0[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[50]),
    .in(in50),
    .out(in_reg_wire_0[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[51]),
    .in(in51),
    .out(in_reg_wire_0[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[52]),
    .in(in52),
    .out(in_reg_wire_0[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[53]),
    .in(in53),
    .out(in_reg_wire_0[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[54]),
    .in(in54),
    .out(in_reg_wire_0[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[55]),
    .in(in55),
    .out(in_reg_wire_0[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[56]),
    .in(in56),
    .out(in_reg_wire_0[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[57]),
    .in(in57),
    .out(in_reg_wire_0[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[58]),
    .in(in58),
    .out(in_reg_wire_0[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[59]),
    .in(in59),
    .out(in_reg_wire_0[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[60]),
    .in(in60),
    .out(in_reg_wire_0[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[61]),
    .in(in61),
    .out(in_reg_wire_0[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[62]),
    .in(in62),
    .out(in_reg_wire_0[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[63]),
    .in(in63),
    .out(in_reg_wire_0[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[64]),
    .in(in64),
    .out(in_reg_wire_0[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[65]),
    .in(in65),
    .out(in_reg_wire_0[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[66]),
    .in(in66),
    .out(in_reg_wire_0[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[67]),
    .in(in67),
    .out(in_reg_wire_0[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[68]),
    .in(in68),
    .out(in_reg_wire_0[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[69]),
    .in(in69),
    .out(in_reg_wire_0[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[70]),
    .in(in70),
    .out(in_reg_wire_0[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[71]),
    .in(in71),
    .out(in_reg_wire_0[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[72]),
    .in(in72),
    .out(in_reg_wire_0[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[73]),
    .in(in73),
    .out(in_reg_wire_0[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[74]),
    .in(in74),
    .out(in_reg_wire_0[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[75]),
    .in(in75),
    .out(in_reg_wire_0[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[76]),
    .in(in76),
    .out(in_reg_wire_0[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[77]),
    .in(in77),
    .out(in_reg_wire_0[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[78]),
    .in(in78),
    .out(in_reg_wire_0[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[79]),
    .in(in79),
    .out(in_reg_wire_0[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[80]),
    .in(in80),
    .out(in_reg_wire_0[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[81]),
    .in(in81),
    .out(in_reg_wire_0[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[82]),
    .in(in82),
    .out(in_reg_wire_0[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[83]),
    .in(in83),
    .out(in_reg_wire_0[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[84]),
    .in(in84),
    .out(in_reg_wire_0[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[85]),
    .in(in85),
    .out(in_reg_wire_0[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[86]),
    .in(in86),
    .out(in_reg_wire_0[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[87]),
    .in(in87),
    .out(in_reg_wire_0[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[88]),
    .in(in88),
    .out(in_reg_wire_0[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[89]),
    .in(in89),
    .out(in_reg_wire_0[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[90]),
    .in(in90),
    .out(in_reg_wire_0[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[91]),
    .in(in91),
    .out(in_reg_wire_0[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[92]),
    .in(in92),
    .out(in_reg_wire_0[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[93]),
    .in(in93),
    .out(in_reg_wire_0[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[94]),
    .in(in94),
    .out(in_reg_wire_0[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[95]),
    .in(in95),
    .out(in_reg_wire_0[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[96]),
    .in(in96),
    .out(in_reg_wire_0[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[97]),
    .in(in97),
    .out(in_reg_wire_0[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[98]),
    .in(in98),
    .out(in_reg_wire_0[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[99]),
    .in(in99),
    .out(in_reg_wire_0[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[100]),
    .in(in100),
    .out(in_reg_wire_0[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[101]),
    .in(in101),
    .out(in_reg_wire_0[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[102]),
    .in(in102),
    .out(in_reg_wire_0[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[103]),
    .in(in103),
    .out(in_reg_wire_0[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[104]),
    .in(in104),
    .out(in_reg_wire_0[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[105]),
    .in(in105),
    .out(in_reg_wire_0[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[106]),
    .in(in106),
    .out(in_reg_wire_0[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[107]),
    .in(in107),
    .out(in_reg_wire_0[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[108]),
    .in(in108),
    .out(in_reg_wire_0[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[109]),
    .in(in109),
    .out(in_reg_wire_0[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[110]),
    .in(in110),
    .out(in_reg_wire_0[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[111]),
    .in(in111),
    .out(in_reg_wire_0[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[112]),
    .in(in112),
    .out(in_reg_wire_0[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[113]),
    .in(in113),
    .out(in_reg_wire_0[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[114]),
    .in(in114),
    .out(in_reg_wire_0[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[115]),
    .in(in115),
    .out(in_reg_wire_0[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[116]),
    .in(in116),
    .out(in_reg_wire_0[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[117]),
    .in(in117),
    .out(in_reg_wire_0[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[118]),
    .in(in118),
    .out(in_reg_wire_0[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[119]),
    .in(in119),
    .out(in_reg_wire_0[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[120]),
    .in(in120),
    .out(in_reg_wire_0[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[121]),
    .in(in121),
    .out(in_reg_wire_0[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[122]),
    .in(in122),
    .out(in_reg_wire_0[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[123]),
    .in(in123),
    .out(in_reg_wire_0[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[124]),
    .in(in124),
    .out(in_reg_wire_0[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[125]),
    .in(in125),
    .out(in_reg_wire_0[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[126]),
    .in(in126),
    .out(in_reg_wire_0[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[127]),
    .in(in127),
    .out(in_reg_wire_0[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[128]),
    .in(in128),
    .out(in_reg_wire_0[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[129]),
    .in(in129),
    .out(in_reg_wire_0[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[130]),
    .in(in130),
    .out(in_reg_wire_0[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[131]),
    .in(in131),
    .out(in_reg_wire_0[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[132]),
    .in(in132),
    .out(in_reg_wire_0[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[133]),
    .in(in133),
    .out(in_reg_wire_0[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[134]),
    .in(in134),
    .out(in_reg_wire_0[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[135]),
    .in(in135),
    .out(in_reg_wire_0[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[136]),
    .in(in136),
    .out(in_reg_wire_0[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[137]),
    .in(in137),
    .out(in_reg_wire_0[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[138]),
    .in(in138),
    .out(in_reg_wire_0[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[139]),
    .in(in139),
    .out(in_reg_wire_0[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[140]),
    .in(in140),
    .out(in_reg_wire_0[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[141]),
    .in(in141),
    .out(in_reg_wire_0[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[142]),
    .in(in142),
    .out(in_reg_wire_0[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[143]),
    .in(in143),
    .out(in_reg_wire_0[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[144]),
    .in(in144),
    .out(in_reg_wire_0[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[145]),
    .in(in145),
    .out(in_reg_wire_0[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[146]),
    .in(in146),
    .out(in_reg_wire_0[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[147]),
    .in(in147),
    .out(in_reg_wire_0[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[148]),
    .in(in148),
    .out(in_reg_wire_0[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[149]),
    .in(in149),
    .out(in_reg_wire_0[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[150]),
    .in(in150),
    .out(in_reg_wire_0[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[151]),
    .in(in151),
    .out(in_reg_wire_0[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[152]),
    .in(in152),
    .out(in_reg_wire_0[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[153]),
    .in(in153),
    .out(in_reg_wire_0[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[154]),
    .in(in154),
    .out(in_reg_wire_0[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[155]),
    .in(in155),
    .out(in_reg_wire_0[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[156]),
    .in(in156),
    .out(in_reg_wire_0[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[157]),
    .in(in157),
    .out(in_reg_wire_0[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[158]),
    .in(in158),
    .out(in_reg_wire_0[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[159]),
    .in(in159),
    .out(in_reg_wire_0[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[160]),
    .in(in160),
    .out(in_reg_wire_0[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[161]),
    .in(in161),
    .out(in_reg_wire_0[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[162]),
    .in(in162),
    .out(in_reg_wire_0[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[163]),
    .in(in163),
    .out(in_reg_wire_0[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[164]),
    .in(in164),
    .out(in_reg_wire_0[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[165]),
    .in(in165),
    .out(in_reg_wire_0[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[166]),
    .in(in166),
    .out(in_reg_wire_0[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[167]),
    .in(in167),
    .out(in_reg_wire_0[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[168]),
    .in(in168),
    .out(in_reg_wire_0[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[169]),
    .in(in169),
    .out(in_reg_wire_0[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[170]),
    .in(in170),
    .out(in_reg_wire_0[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[171]),
    .in(in171),
    .out(in_reg_wire_0[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[172]),
    .in(in172),
    .out(in_reg_wire_0[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[173]),
    .in(in173),
    .out(in_reg_wire_0[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[174]),
    .in(in174),
    .out(in_reg_wire_0[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[175]),
    .in(in175),
    .out(in_reg_wire_0[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[176]),
    .in(in176),
    .out(in_reg_wire_0[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[177]),
    .in(in177),
    .out(in_reg_wire_0[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[178]),
    .in(in178),
    .out(in_reg_wire_0[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[179]),
    .in(in179),
    .out(in_reg_wire_0[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[180]),
    .in(in180),
    .out(in_reg_wire_0[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[181]),
    .in(in181),
    .out(in_reg_wire_0[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[182]),
    .in(in182),
    .out(in_reg_wire_0[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[183]),
    .in(in183),
    .out(in_reg_wire_0[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[184]),
    .in(in184),
    .out(in_reg_wire_0[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[185]),
    .in(in185),
    .out(in_reg_wire_0[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[186]),
    .in(in186),
    .out(in_reg_wire_0[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[187]),
    .in(in187),
    .out(in_reg_wire_0[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[188]),
    .in(in188),
    .out(in_reg_wire_0[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[189]),
    .in(in189),
    .out(in_reg_wire_0[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[190]),
    .in(in190),
    .out(in_reg_wire_0[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[191]),
    .in(in191),
    .out(in_reg_wire_0[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[192]),
    .in(in192),
    .out(in_reg_wire_0[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[193]),
    .in(in193),
    .out(in_reg_wire_0[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[194]),
    .in(in194),
    .out(in_reg_wire_0[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[195]),
    .in(in195),
    .out(in_reg_wire_0[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[196]),
    .in(in196),
    .out(in_reg_wire_0[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[197]),
    .in(in197),
    .out(in_reg_wire_0[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[198]),
    .in(in198),
    .out(in_reg_wire_0[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[199]),
    .in(in199),
    .out(in_reg_wire_0[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[200]),
    .in(in200),
    .out(in_reg_wire_0[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[201]),
    .in(in201),
    .out(in_reg_wire_0[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[202]),
    .in(in202),
    .out(in_reg_wire_0[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[203]),
    .in(in203),
    .out(in_reg_wire_0[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[204]),
    .in(in204),
    .out(in_reg_wire_0[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[205]),
    .in(in205),
    .out(in_reg_wire_0[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[206]),
    .in(in206),
    .out(in_reg_wire_0[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[207]),
    .in(in207),
    .out(in_reg_wire_0[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[208]),
    .in(in208),
    .out(in_reg_wire_0[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[209]),
    .in(in209),
    .out(in_reg_wire_0[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[210]),
    .in(in210),
    .out(in_reg_wire_0[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[211]),
    .in(in211),
    .out(in_reg_wire_0[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[212]),
    .in(in212),
    .out(in_reg_wire_0[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[213]),
    .in(in213),
    .out(in_reg_wire_0[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[214]),
    .in(in214),
    .out(in_reg_wire_0[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[215]),
    .in(in215),
    .out(in_reg_wire_0[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[216]),
    .in(in216),
    .out(in_reg_wire_0[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[217]),
    .in(in217),
    .out(in_reg_wire_0[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[218]),
    .in(in218),
    .out(in_reg_wire_0[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[219]),
    .in(in219),
    .out(in_reg_wire_0[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[220]),
    .in(in220),
    .out(in_reg_wire_0[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[221]),
    .in(in221),
    .out(in_reg_wire_0[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[222]),
    .in(in222),
    .out(in_reg_wire_0[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[223]),
    .in(in223),
    .out(in_reg_wire_0[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[224]),
    .in(in224),
    .out(in_reg_wire_0[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[225]),
    .in(in225),
    .out(in_reg_wire_0[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[226]),
    .in(in226),
    .out(in_reg_wire_0[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[227]),
    .in(in227),
    .out(in_reg_wire_0[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[228]),
    .in(in228),
    .out(in_reg_wire_0[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[229]),
    .in(in229),
    .out(in_reg_wire_0[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[230]),
    .in(in230),
    .out(in_reg_wire_0[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[231]),
    .in(in231),
    .out(in_reg_wire_0[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[232]),
    .in(in232),
    .out(in_reg_wire_0[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[233]),
    .in(in233),
    .out(in_reg_wire_0[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[234]),
    .in(in234),
    .out(in_reg_wire_0[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[235]),
    .in(in235),
    .out(in_reg_wire_0[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[236]),
    .in(in236),
    .out(in_reg_wire_0[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[237]),
    .in(in237),
    .out(in_reg_wire_0[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[238]),
    .in(in238),
    .out(in_reg_wire_0[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[239]),
    .in(in239),
    .out(in_reg_wire_0[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[240]),
    .in(in240),
    .out(in_reg_wire_0[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[241]),
    .in(in241),
    .out(in_reg_wire_0[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[242]),
    .in(in242),
    .out(in_reg_wire_0[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[243]),
    .in(in243),
    .out(in_reg_wire_0[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[244]),
    .in(in244),
    .out(in_reg_wire_0[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[245]),
    .in(in245),
    .out(in_reg_wire_0[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[246]),
    .in(in246),
    .out(in_reg_wire_0[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[247]),
    .in(in247),
    .out(in_reg_wire_0[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[248]),
    .in(in248),
    .out(in_reg_wire_0[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[249]),
    .in(in249),
    .out(in_reg_wire_0[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[250]),
    .in(in250),
    .out(in_reg_wire_0[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[251]),
    .in(in251),
    .out(in_reg_wire_0[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[252]),
    .in(in252),
    .out(in_reg_wire_0[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[253]),
    .in(in253),
    .out(in_reg_wire_0[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[254]),
    .in(in254),
    .out(in_reg_wire_0[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[255]),
    .in(in255),
    .out(in_reg_wire_0[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[256]),
    .in(in_reg_wire_1[0]),
    .out(in_reg_wire_2[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[257]),
    .in(in_reg_wire_1[1]),
    .out(in_reg_wire_2[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[258]),
    .in(in_reg_wire_1[2]),
    .out(in_reg_wire_2[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[259]),
    .in(in_reg_wire_1[3]),
    .out(in_reg_wire_2[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[260]),
    .in(in_reg_wire_1[4]),
    .out(in_reg_wire_2[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[261]),
    .in(in_reg_wire_1[5]),
    .out(in_reg_wire_2[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[262]),
    .in(in_reg_wire_1[6]),
    .out(in_reg_wire_2[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[263]),
    .in(in_reg_wire_1[7]),
    .out(in_reg_wire_2[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[264]),
    .in(in_reg_wire_1[8]),
    .out(in_reg_wire_2[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[265]),
    .in(in_reg_wire_1[9]),
    .out(in_reg_wire_2[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[266]),
    .in(in_reg_wire_1[10]),
    .out(in_reg_wire_2[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[267]),
    .in(in_reg_wire_1[11]),
    .out(in_reg_wire_2[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[268]),
    .in(in_reg_wire_1[12]),
    .out(in_reg_wire_2[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[269]),
    .in(in_reg_wire_1[13]),
    .out(in_reg_wire_2[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[270]),
    .in(in_reg_wire_1[14]),
    .out(in_reg_wire_2[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[271]),
    .in(in_reg_wire_1[15]),
    .out(in_reg_wire_2[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[272]),
    .in(in_reg_wire_1[16]),
    .out(in_reg_wire_2[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[273]),
    .in(in_reg_wire_1[17]),
    .out(in_reg_wire_2[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[274]),
    .in(in_reg_wire_1[18]),
    .out(in_reg_wire_2[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[275]),
    .in(in_reg_wire_1[19]),
    .out(in_reg_wire_2[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[276]),
    .in(in_reg_wire_1[20]),
    .out(in_reg_wire_2[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[277]),
    .in(in_reg_wire_1[21]),
    .out(in_reg_wire_2[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[278]),
    .in(in_reg_wire_1[22]),
    .out(in_reg_wire_2[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[279]),
    .in(in_reg_wire_1[23]),
    .out(in_reg_wire_2[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[280]),
    .in(in_reg_wire_1[24]),
    .out(in_reg_wire_2[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[281]),
    .in(in_reg_wire_1[25]),
    .out(in_reg_wire_2[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[282]),
    .in(in_reg_wire_1[26]),
    .out(in_reg_wire_2[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[283]),
    .in(in_reg_wire_1[27]),
    .out(in_reg_wire_2[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[284]),
    .in(in_reg_wire_1[28]),
    .out(in_reg_wire_2[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[285]),
    .in(in_reg_wire_1[29]),
    .out(in_reg_wire_2[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[286]),
    .in(in_reg_wire_1[30]),
    .out(in_reg_wire_2[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[287]),
    .in(in_reg_wire_1[31]),
    .out(in_reg_wire_2[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[288]),
    .in(in_reg_wire_1[32]),
    .out(in_reg_wire_2[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[289]),
    .in(in_reg_wire_1[33]),
    .out(in_reg_wire_2[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[290]),
    .in(in_reg_wire_1[34]),
    .out(in_reg_wire_2[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[291]),
    .in(in_reg_wire_1[35]),
    .out(in_reg_wire_2[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[292]),
    .in(in_reg_wire_1[36]),
    .out(in_reg_wire_2[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[293]),
    .in(in_reg_wire_1[37]),
    .out(in_reg_wire_2[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[294]),
    .in(in_reg_wire_1[38]),
    .out(in_reg_wire_2[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[295]),
    .in(in_reg_wire_1[39]),
    .out(in_reg_wire_2[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[296]),
    .in(in_reg_wire_1[40]),
    .out(in_reg_wire_2[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[297]),
    .in(in_reg_wire_1[41]),
    .out(in_reg_wire_2[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[298]),
    .in(in_reg_wire_1[42]),
    .out(in_reg_wire_2[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[299]),
    .in(in_reg_wire_1[43]),
    .out(in_reg_wire_2[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[300]),
    .in(in_reg_wire_1[44]),
    .out(in_reg_wire_2[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[301]),
    .in(in_reg_wire_1[45]),
    .out(in_reg_wire_2[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[302]),
    .in(in_reg_wire_1[46]),
    .out(in_reg_wire_2[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[303]),
    .in(in_reg_wire_1[47]),
    .out(in_reg_wire_2[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[304]),
    .in(in_reg_wire_1[48]),
    .out(in_reg_wire_2[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[305]),
    .in(in_reg_wire_1[49]),
    .out(in_reg_wire_2[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[306]),
    .in(in_reg_wire_1[50]),
    .out(in_reg_wire_2[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[307]),
    .in(in_reg_wire_1[51]),
    .out(in_reg_wire_2[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[308]),
    .in(in_reg_wire_1[52]),
    .out(in_reg_wire_2[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[309]),
    .in(in_reg_wire_1[53]),
    .out(in_reg_wire_2[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[310]),
    .in(in_reg_wire_1[54]),
    .out(in_reg_wire_2[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[311]),
    .in(in_reg_wire_1[55]),
    .out(in_reg_wire_2[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[312]),
    .in(in_reg_wire_1[56]),
    .out(in_reg_wire_2[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[313]),
    .in(in_reg_wire_1[57]),
    .out(in_reg_wire_2[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[314]),
    .in(in_reg_wire_1[58]),
    .out(in_reg_wire_2[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[315]),
    .in(in_reg_wire_1[59]),
    .out(in_reg_wire_2[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[316]),
    .in(in_reg_wire_1[60]),
    .out(in_reg_wire_2[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[317]),
    .in(in_reg_wire_1[61]),
    .out(in_reg_wire_2[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[318]),
    .in(in_reg_wire_1[62]),
    .out(in_reg_wire_2[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[319]),
    .in(in_reg_wire_1[63]),
    .out(in_reg_wire_2[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[320]),
    .in(in_reg_wire_1[64]),
    .out(in_reg_wire_2[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[321]),
    .in(in_reg_wire_1[65]),
    .out(in_reg_wire_2[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[322]),
    .in(in_reg_wire_1[66]),
    .out(in_reg_wire_2[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[323]),
    .in(in_reg_wire_1[67]),
    .out(in_reg_wire_2[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[324]),
    .in(in_reg_wire_1[68]),
    .out(in_reg_wire_2[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[325]),
    .in(in_reg_wire_1[69]),
    .out(in_reg_wire_2[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[326]),
    .in(in_reg_wire_1[70]),
    .out(in_reg_wire_2[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[327]),
    .in(in_reg_wire_1[71]),
    .out(in_reg_wire_2[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[328]),
    .in(in_reg_wire_1[72]),
    .out(in_reg_wire_2[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[329]),
    .in(in_reg_wire_1[73]),
    .out(in_reg_wire_2[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[330]),
    .in(in_reg_wire_1[74]),
    .out(in_reg_wire_2[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[331]),
    .in(in_reg_wire_1[75]),
    .out(in_reg_wire_2[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[332]),
    .in(in_reg_wire_1[76]),
    .out(in_reg_wire_2[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[333]),
    .in(in_reg_wire_1[77]),
    .out(in_reg_wire_2[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[334]),
    .in(in_reg_wire_1[78]),
    .out(in_reg_wire_2[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[335]),
    .in(in_reg_wire_1[79]),
    .out(in_reg_wire_2[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[336]),
    .in(in_reg_wire_1[80]),
    .out(in_reg_wire_2[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[337]),
    .in(in_reg_wire_1[81]),
    .out(in_reg_wire_2[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[338]),
    .in(in_reg_wire_1[82]),
    .out(in_reg_wire_2[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[339]),
    .in(in_reg_wire_1[83]),
    .out(in_reg_wire_2[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[340]),
    .in(in_reg_wire_1[84]),
    .out(in_reg_wire_2[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[341]),
    .in(in_reg_wire_1[85]),
    .out(in_reg_wire_2[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[342]),
    .in(in_reg_wire_1[86]),
    .out(in_reg_wire_2[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[343]),
    .in(in_reg_wire_1[87]),
    .out(in_reg_wire_2[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[344]),
    .in(in_reg_wire_1[88]),
    .out(in_reg_wire_2[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[345]),
    .in(in_reg_wire_1[89]),
    .out(in_reg_wire_2[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[346]),
    .in(in_reg_wire_1[90]),
    .out(in_reg_wire_2[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[347]),
    .in(in_reg_wire_1[91]),
    .out(in_reg_wire_2[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[348]),
    .in(in_reg_wire_1[92]),
    .out(in_reg_wire_2[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[349]),
    .in(in_reg_wire_1[93]),
    .out(in_reg_wire_2[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[350]),
    .in(in_reg_wire_1[94]),
    .out(in_reg_wire_2[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[351]),
    .in(in_reg_wire_1[95]),
    .out(in_reg_wire_2[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[352]),
    .in(in_reg_wire_1[96]),
    .out(in_reg_wire_2[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[353]),
    .in(in_reg_wire_1[97]),
    .out(in_reg_wire_2[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[354]),
    .in(in_reg_wire_1[98]),
    .out(in_reg_wire_2[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[355]),
    .in(in_reg_wire_1[99]),
    .out(in_reg_wire_2[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[356]),
    .in(in_reg_wire_1[100]),
    .out(in_reg_wire_2[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[357]),
    .in(in_reg_wire_1[101]),
    .out(in_reg_wire_2[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[358]),
    .in(in_reg_wire_1[102]),
    .out(in_reg_wire_2[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[359]),
    .in(in_reg_wire_1[103]),
    .out(in_reg_wire_2[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[360]),
    .in(in_reg_wire_1[104]),
    .out(in_reg_wire_2[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[361]),
    .in(in_reg_wire_1[105]),
    .out(in_reg_wire_2[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[362]),
    .in(in_reg_wire_1[106]),
    .out(in_reg_wire_2[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[363]),
    .in(in_reg_wire_1[107]),
    .out(in_reg_wire_2[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[364]),
    .in(in_reg_wire_1[108]),
    .out(in_reg_wire_2[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[365]),
    .in(in_reg_wire_1[109]),
    .out(in_reg_wire_2[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[366]),
    .in(in_reg_wire_1[110]),
    .out(in_reg_wire_2[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[367]),
    .in(in_reg_wire_1[111]),
    .out(in_reg_wire_2[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[368]),
    .in(in_reg_wire_1[112]),
    .out(in_reg_wire_2[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[369]),
    .in(in_reg_wire_1[113]),
    .out(in_reg_wire_2[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[370]),
    .in(in_reg_wire_1[114]),
    .out(in_reg_wire_2[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[371]),
    .in(in_reg_wire_1[115]),
    .out(in_reg_wire_2[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[372]),
    .in(in_reg_wire_1[116]),
    .out(in_reg_wire_2[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[373]),
    .in(in_reg_wire_1[117]),
    .out(in_reg_wire_2[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[374]),
    .in(in_reg_wire_1[118]),
    .out(in_reg_wire_2[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[375]),
    .in(in_reg_wire_1[119]),
    .out(in_reg_wire_2[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[376]),
    .in(in_reg_wire_1[120]),
    .out(in_reg_wire_2[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[377]),
    .in(in_reg_wire_1[121]),
    .out(in_reg_wire_2[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[378]),
    .in(in_reg_wire_1[122]),
    .out(in_reg_wire_2[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[379]),
    .in(in_reg_wire_1[123]),
    .out(in_reg_wire_2[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[380]),
    .in(in_reg_wire_1[124]),
    .out(in_reg_wire_2[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[381]),
    .in(in_reg_wire_1[125]),
    .out(in_reg_wire_2[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[382]),
    .in(in_reg_wire_1[126]),
    .out(in_reg_wire_2[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[383]),
    .in(in_reg_wire_1[127]),
    .out(in_reg_wire_2[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[384]),
    .in(in_reg_wire_1[128]),
    .out(in_reg_wire_2[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[385]),
    .in(in_reg_wire_1[129]),
    .out(in_reg_wire_2[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[386]),
    .in(in_reg_wire_1[130]),
    .out(in_reg_wire_2[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[387]),
    .in(in_reg_wire_1[131]),
    .out(in_reg_wire_2[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[388]),
    .in(in_reg_wire_1[132]),
    .out(in_reg_wire_2[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[389]),
    .in(in_reg_wire_1[133]),
    .out(in_reg_wire_2[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[390]),
    .in(in_reg_wire_1[134]),
    .out(in_reg_wire_2[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[391]),
    .in(in_reg_wire_1[135]),
    .out(in_reg_wire_2[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[392]),
    .in(in_reg_wire_1[136]),
    .out(in_reg_wire_2[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[393]),
    .in(in_reg_wire_1[137]),
    .out(in_reg_wire_2[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[394]),
    .in(in_reg_wire_1[138]),
    .out(in_reg_wire_2[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[395]),
    .in(in_reg_wire_1[139]),
    .out(in_reg_wire_2[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[396]),
    .in(in_reg_wire_1[140]),
    .out(in_reg_wire_2[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[397]),
    .in(in_reg_wire_1[141]),
    .out(in_reg_wire_2[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[398]),
    .in(in_reg_wire_1[142]),
    .out(in_reg_wire_2[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[399]),
    .in(in_reg_wire_1[143]),
    .out(in_reg_wire_2[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[400]),
    .in(in_reg_wire_1[144]),
    .out(in_reg_wire_2[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[401]),
    .in(in_reg_wire_1[145]),
    .out(in_reg_wire_2[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[402]),
    .in(in_reg_wire_1[146]),
    .out(in_reg_wire_2[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[403]),
    .in(in_reg_wire_1[147]),
    .out(in_reg_wire_2[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[404]),
    .in(in_reg_wire_1[148]),
    .out(in_reg_wire_2[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[405]),
    .in(in_reg_wire_1[149]),
    .out(in_reg_wire_2[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[406]),
    .in(in_reg_wire_1[150]),
    .out(in_reg_wire_2[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[407]),
    .in(in_reg_wire_1[151]),
    .out(in_reg_wire_2[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[408]),
    .in(in_reg_wire_1[152]),
    .out(in_reg_wire_2[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[409]),
    .in(in_reg_wire_1[153]),
    .out(in_reg_wire_2[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[410]),
    .in(in_reg_wire_1[154]),
    .out(in_reg_wire_2[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[411]),
    .in(in_reg_wire_1[155]),
    .out(in_reg_wire_2[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[412]),
    .in(in_reg_wire_1[156]),
    .out(in_reg_wire_2[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[413]),
    .in(in_reg_wire_1[157]),
    .out(in_reg_wire_2[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[414]),
    .in(in_reg_wire_1[158]),
    .out(in_reg_wire_2[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[415]),
    .in(in_reg_wire_1[159]),
    .out(in_reg_wire_2[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[416]),
    .in(in_reg_wire_1[160]),
    .out(in_reg_wire_2[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[417]),
    .in(in_reg_wire_1[161]),
    .out(in_reg_wire_2[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[418]),
    .in(in_reg_wire_1[162]),
    .out(in_reg_wire_2[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[419]),
    .in(in_reg_wire_1[163]),
    .out(in_reg_wire_2[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[420]),
    .in(in_reg_wire_1[164]),
    .out(in_reg_wire_2[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[421]),
    .in(in_reg_wire_1[165]),
    .out(in_reg_wire_2[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[422]),
    .in(in_reg_wire_1[166]),
    .out(in_reg_wire_2[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[423]),
    .in(in_reg_wire_1[167]),
    .out(in_reg_wire_2[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[424]),
    .in(in_reg_wire_1[168]),
    .out(in_reg_wire_2[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[425]),
    .in(in_reg_wire_1[169]),
    .out(in_reg_wire_2[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[426]),
    .in(in_reg_wire_1[170]),
    .out(in_reg_wire_2[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[427]),
    .in(in_reg_wire_1[171]),
    .out(in_reg_wire_2[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[428]),
    .in(in_reg_wire_1[172]),
    .out(in_reg_wire_2[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[429]),
    .in(in_reg_wire_1[173]),
    .out(in_reg_wire_2[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[430]),
    .in(in_reg_wire_1[174]),
    .out(in_reg_wire_2[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[431]),
    .in(in_reg_wire_1[175]),
    .out(in_reg_wire_2[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[432]),
    .in(in_reg_wire_1[176]),
    .out(in_reg_wire_2[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[433]),
    .in(in_reg_wire_1[177]),
    .out(in_reg_wire_2[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[434]),
    .in(in_reg_wire_1[178]),
    .out(in_reg_wire_2[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[435]),
    .in(in_reg_wire_1[179]),
    .out(in_reg_wire_2[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[436]),
    .in(in_reg_wire_1[180]),
    .out(in_reg_wire_2[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[437]),
    .in(in_reg_wire_1[181]),
    .out(in_reg_wire_2[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[438]),
    .in(in_reg_wire_1[182]),
    .out(in_reg_wire_2[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[439]),
    .in(in_reg_wire_1[183]),
    .out(in_reg_wire_2[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[440]),
    .in(in_reg_wire_1[184]),
    .out(in_reg_wire_2[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[441]),
    .in(in_reg_wire_1[185]),
    .out(in_reg_wire_2[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[442]),
    .in(in_reg_wire_1[186]),
    .out(in_reg_wire_2[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[443]),
    .in(in_reg_wire_1[187]),
    .out(in_reg_wire_2[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[444]),
    .in(in_reg_wire_1[188]),
    .out(in_reg_wire_2[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[445]),
    .in(in_reg_wire_1[189]),
    .out(in_reg_wire_2[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[446]),
    .in(in_reg_wire_1[190]),
    .out(in_reg_wire_2[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[447]),
    .in(in_reg_wire_1[191]),
    .out(in_reg_wire_2[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[448]),
    .in(in_reg_wire_1[192]),
    .out(in_reg_wire_2[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[449]),
    .in(in_reg_wire_1[193]),
    .out(in_reg_wire_2[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[450]),
    .in(in_reg_wire_1[194]),
    .out(in_reg_wire_2[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[451]),
    .in(in_reg_wire_1[195]),
    .out(in_reg_wire_2[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[452]),
    .in(in_reg_wire_1[196]),
    .out(in_reg_wire_2[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[453]),
    .in(in_reg_wire_1[197]),
    .out(in_reg_wire_2[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[454]),
    .in(in_reg_wire_1[198]),
    .out(in_reg_wire_2[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[455]),
    .in(in_reg_wire_1[199]),
    .out(in_reg_wire_2[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[456]),
    .in(in_reg_wire_1[200]),
    .out(in_reg_wire_2[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[457]),
    .in(in_reg_wire_1[201]),
    .out(in_reg_wire_2[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[458]),
    .in(in_reg_wire_1[202]),
    .out(in_reg_wire_2[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[459]),
    .in(in_reg_wire_1[203]),
    .out(in_reg_wire_2[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[460]),
    .in(in_reg_wire_1[204]),
    .out(in_reg_wire_2[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[461]),
    .in(in_reg_wire_1[205]),
    .out(in_reg_wire_2[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[462]),
    .in(in_reg_wire_1[206]),
    .out(in_reg_wire_2[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[463]),
    .in(in_reg_wire_1[207]),
    .out(in_reg_wire_2[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[464]),
    .in(in_reg_wire_1[208]),
    .out(in_reg_wire_2[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[465]),
    .in(in_reg_wire_1[209]),
    .out(in_reg_wire_2[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[466]),
    .in(in_reg_wire_1[210]),
    .out(in_reg_wire_2[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[467]),
    .in(in_reg_wire_1[211]),
    .out(in_reg_wire_2[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[468]),
    .in(in_reg_wire_1[212]),
    .out(in_reg_wire_2[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[469]),
    .in(in_reg_wire_1[213]),
    .out(in_reg_wire_2[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[470]),
    .in(in_reg_wire_1[214]),
    .out(in_reg_wire_2[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[471]),
    .in(in_reg_wire_1[215]),
    .out(in_reg_wire_2[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[472]),
    .in(in_reg_wire_1[216]),
    .out(in_reg_wire_2[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[473]),
    .in(in_reg_wire_1[217]),
    .out(in_reg_wire_2[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[474]),
    .in(in_reg_wire_1[218]),
    .out(in_reg_wire_2[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[475]),
    .in(in_reg_wire_1[219]),
    .out(in_reg_wire_2[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[476]),
    .in(in_reg_wire_1[220]),
    .out(in_reg_wire_2[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[477]),
    .in(in_reg_wire_1[221]),
    .out(in_reg_wire_2[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[478]),
    .in(in_reg_wire_1[222]),
    .out(in_reg_wire_2[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[479]),
    .in(in_reg_wire_1[223]),
    .out(in_reg_wire_2[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[480]),
    .in(in_reg_wire_1[224]),
    .out(in_reg_wire_2[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[481]),
    .in(in_reg_wire_1[225]),
    .out(in_reg_wire_2[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[482]),
    .in(in_reg_wire_1[226]),
    .out(in_reg_wire_2[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[483]),
    .in(in_reg_wire_1[227]),
    .out(in_reg_wire_2[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[484]),
    .in(in_reg_wire_1[228]),
    .out(in_reg_wire_2[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[485]),
    .in(in_reg_wire_1[229]),
    .out(in_reg_wire_2[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[486]),
    .in(in_reg_wire_1[230]),
    .out(in_reg_wire_2[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[487]),
    .in(in_reg_wire_1[231]),
    .out(in_reg_wire_2[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[488]),
    .in(in_reg_wire_1[232]),
    .out(in_reg_wire_2[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[489]),
    .in(in_reg_wire_1[233]),
    .out(in_reg_wire_2[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[490]),
    .in(in_reg_wire_1[234]),
    .out(in_reg_wire_2[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[491]),
    .in(in_reg_wire_1[235]),
    .out(in_reg_wire_2[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[492]),
    .in(in_reg_wire_1[236]),
    .out(in_reg_wire_2[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[493]),
    .in(in_reg_wire_1[237]),
    .out(in_reg_wire_2[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[494]),
    .in(in_reg_wire_1[238]),
    .out(in_reg_wire_2[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[495]),
    .in(in_reg_wire_1[239]),
    .out(in_reg_wire_2[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[496]),
    .in(in_reg_wire_1[240]),
    .out(in_reg_wire_2[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[497]),
    .in(in_reg_wire_1[241]),
    .out(in_reg_wire_2[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[498]),
    .in(in_reg_wire_1[242]),
    .out(in_reg_wire_2[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[499]),
    .in(in_reg_wire_1[243]),
    .out(in_reg_wire_2[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[500]),
    .in(in_reg_wire_1[244]),
    .out(in_reg_wire_2[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[501]),
    .in(in_reg_wire_1[245]),
    .out(in_reg_wire_2[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[502]),
    .in(in_reg_wire_1[246]),
    .out(in_reg_wire_2[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[503]),
    .in(in_reg_wire_1[247]),
    .out(in_reg_wire_2[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[504]),
    .in(in_reg_wire_1[248]),
    .out(in_reg_wire_2[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[505]),
    .in(in_reg_wire_1[249]),
    .out(in_reg_wire_2[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[506]),
    .in(in_reg_wire_1[250]),
    .out(in_reg_wire_2[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[507]),
    .in(in_reg_wire_1[251]),
    .out(in_reg_wire_2[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[508]),
    .in(in_reg_wire_1[252]),
    .out(in_reg_wire_2[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[509]),
    .in(in_reg_wire_1[253]),
    .out(in_reg_wire_2[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[510]),
    .in(in_reg_wire_1[254]),
    .out(in_reg_wire_2[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[511]),
    .in(in_reg_wire_1[255]),
    .out(in_reg_wire_2[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[512]),
    .in(in_reg_wire_3[0]),
    .out(in_reg_wire_4[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[513]),
    .in(in_reg_wire_3[1]),
    .out(in_reg_wire_4[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[514]),
    .in(in_reg_wire_3[2]),
    .out(in_reg_wire_4[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[515]),
    .in(in_reg_wire_3[3]),
    .out(in_reg_wire_4[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[516]),
    .in(in_reg_wire_3[4]),
    .out(in_reg_wire_4[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[517]),
    .in(in_reg_wire_3[5]),
    .out(in_reg_wire_4[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[518]),
    .in(in_reg_wire_3[6]),
    .out(in_reg_wire_4[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[519]),
    .in(in_reg_wire_3[7]),
    .out(in_reg_wire_4[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[520]),
    .in(in_reg_wire_3[8]),
    .out(in_reg_wire_4[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[521]),
    .in(in_reg_wire_3[9]),
    .out(in_reg_wire_4[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[522]),
    .in(in_reg_wire_3[10]),
    .out(in_reg_wire_4[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[523]),
    .in(in_reg_wire_3[11]),
    .out(in_reg_wire_4[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[524]),
    .in(in_reg_wire_3[12]),
    .out(in_reg_wire_4[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[525]),
    .in(in_reg_wire_3[13]),
    .out(in_reg_wire_4[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[526]),
    .in(in_reg_wire_3[14]),
    .out(in_reg_wire_4[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[527]),
    .in(in_reg_wire_3[15]),
    .out(in_reg_wire_4[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[528]),
    .in(in_reg_wire_3[16]),
    .out(in_reg_wire_4[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[529]),
    .in(in_reg_wire_3[17]),
    .out(in_reg_wire_4[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[530]),
    .in(in_reg_wire_3[18]),
    .out(in_reg_wire_4[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[531]),
    .in(in_reg_wire_3[19]),
    .out(in_reg_wire_4[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[532]),
    .in(in_reg_wire_3[20]),
    .out(in_reg_wire_4[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[533]),
    .in(in_reg_wire_3[21]),
    .out(in_reg_wire_4[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[534]),
    .in(in_reg_wire_3[22]),
    .out(in_reg_wire_4[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[535]),
    .in(in_reg_wire_3[23]),
    .out(in_reg_wire_4[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[536]),
    .in(in_reg_wire_3[24]),
    .out(in_reg_wire_4[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[537]),
    .in(in_reg_wire_3[25]),
    .out(in_reg_wire_4[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[538]),
    .in(in_reg_wire_3[26]),
    .out(in_reg_wire_4[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[539]),
    .in(in_reg_wire_3[27]),
    .out(in_reg_wire_4[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[540]),
    .in(in_reg_wire_3[28]),
    .out(in_reg_wire_4[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[541]),
    .in(in_reg_wire_3[29]),
    .out(in_reg_wire_4[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[542]),
    .in(in_reg_wire_3[30]),
    .out(in_reg_wire_4[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[543]),
    .in(in_reg_wire_3[31]),
    .out(in_reg_wire_4[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[544]),
    .in(in_reg_wire_3[32]),
    .out(in_reg_wire_4[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[545]),
    .in(in_reg_wire_3[33]),
    .out(in_reg_wire_4[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[546]),
    .in(in_reg_wire_3[34]),
    .out(in_reg_wire_4[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[547]),
    .in(in_reg_wire_3[35]),
    .out(in_reg_wire_4[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[548]),
    .in(in_reg_wire_3[36]),
    .out(in_reg_wire_4[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[549]),
    .in(in_reg_wire_3[37]),
    .out(in_reg_wire_4[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[550]),
    .in(in_reg_wire_3[38]),
    .out(in_reg_wire_4[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[551]),
    .in(in_reg_wire_3[39]),
    .out(in_reg_wire_4[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[552]),
    .in(in_reg_wire_3[40]),
    .out(in_reg_wire_4[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[553]),
    .in(in_reg_wire_3[41]),
    .out(in_reg_wire_4[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[554]),
    .in(in_reg_wire_3[42]),
    .out(in_reg_wire_4[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[555]),
    .in(in_reg_wire_3[43]),
    .out(in_reg_wire_4[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[556]),
    .in(in_reg_wire_3[44]),
    .out(in_reg_wire_4[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[557]),
    .in(in_reg_wire_3[45]),
    .out(in_reg_wire_4[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[558]),
    .in(in_reg_wire_3[46]),
    .out(in_reg_wire_4[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[559]),
    .in(in_reg_wire_3[47]),
    .out(in_reg_wire_4[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[560]),
    .in(in_reg_wire_3[48]),
    .out(in_reg_wire_4[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[561]),
    .in(in_reg_wire_3[49]),
    .out(in_reg_wire_4[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[562]),
    .in(in_reg_wire_3[50]),
    .out(in_reg_wire_4[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[563]),
    .in(in_reg_wire_3[51]),
    .out(in_reg_wire_4[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[564]),
    .in(in_reg_wire_3[52]),
    .out(in_reg_wire_4[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[565]),
    .in(in_reg_wire_3[53]),
    .out(in_reg_wire_4[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[566]),
    .in(in_reg_wire_3[54]),
    .out(in_reg_wire_4[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[567]),
    .in(in_reg_wire_3[55]),
    .out(in_reg_wire_4[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[568]),
    .in(in_reg_wire_3[56]),
    .out(in_reg_wire_4[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[569]),
    .in(in_reg_wire_3[57]),
    .out(in_reg_wire_4[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[570]),
    .in(in_reg_wire_3[58]),
    .out(in_reg_wire_4[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[571]),
    .in(in_reg_wire_3[59]),
    .out(in_reg_wire_4[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[572]),
    .in(in_reg_wire_3[60]),
    .out(in_reg_wire_4[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[573]),
    .in(in_reg_wire_3[61]),
    .out(in_reg_wire_4[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[574]),
    .in(in_reg_wire_3[62]),
    .out(in_reg_wire_4[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[575]),
    .in(in_reg_wire_3[63]),
    .out(in_reg_wire_4[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[576]),
    .in(in_reg_wire_3[64]),
    .out(in_reg_wire_4[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[577]),
    .in(in_reg_wire_3[65]),
    .out(in_reg_wire_4[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[578]),
    .in(in_reg_wire_3[66]),
    .out(in_reg_wire_4[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[579]),
    .in(in_reg_wire_3[67]),
    .out(in_reg_wire_4[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[580]),
    .in(in_reg_wire_3[68]),
    .out(in_reg_wire_4[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[581]),
    .in(in_reg_wire_3[69]),
    .out(in_reg_wire_4[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[582]),
    .in(in_reg_wire_3[70]),
    .out(in_reg_wire_4[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[583]),
    .in(in_reg_wire_3[71]),
    .out(in_reg_wire_4[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[584]),
    .in(in_reg_wire_3[72]),
    .out(in_reg_wire_4[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[585]),
    .in(in_reg_wire_3[73]),
    .out(in_reg_wire_4[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[586]),
    .in(in_reg_wire_3[74]),
    .out(in_reg_wire_4[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[587]),
    .in(in_reg_wire_3[75]),
    .out(in_reg_wire_4[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[588]),
    .in(in_reg_wire_3[76]),
    .out(in_reg_wire_4[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[589]),
    .in(in_reg_wire_3[77]),
    .out(in_reg_wire_4[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[590]),
    .in(in_reg_wire_3[78]),
    .out(in_reg_wire_4[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[591]),
    .in(in_reg_wire_3[79]),
    .out(in_reg_wire_4[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[592]),
    .in(in_reg_wire_3[80]),
    .out(in_reg_wire_4[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[593]),
    .in(in_reg_wire_3[81]),
    .out(in_reg_wire_4[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[594]),
    .in(in_reg_wire_3[82]),
    .out(in_reg_wire_4[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[595]),
    .in(in_reg_wire_3[83]),
    .out(in_reg_wire_4[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[596]),
    .in(in_reg_wire_3[84]),
    .out(in_reg_wire_4[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[597]),
    .in(in_reg_wire_3[85]),
    .out(in_reg_wire_4[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[598]),
    .in(in_reg_wire_3[86]),
    .out(in_reg_wire_4[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[599]),
    .in(in_reg_wire_3[87]),
    .out(in_reg_wire_4[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[600]),
    .in(in_reg_wire_3[88]),
    .out(in_reg_wire_4[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[601]),
    .in(in_reg_wire_3[89]),
    .out(in_reg_wire_4[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[602]),
    .in(in_reg_wire_3[90]),
    .out(in_reg_wire_4[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[603]),
    .in(in_reg_wire_3[91]),
    .out(in_reg_wire_4[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[604]),
    .in(in_reg_wire_3[92]),
    .out(in_reg_wire_4[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[605]),
    .in(in_reg_wire_3[93]),
    .out(in_reg_wire_4[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[606]),
    .in(in_reg_wire_3[94]),
    .out(in_reg_wire_4[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[607]),
    .in(in_reg_wire_3[95]),
    .out(in_reg_wire_4[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[608]),
    .in(in_reg_wire_3[96]),
    .out(in_reg_wire_4[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[609]),
    .in(in_reg_wire_3[97]),
    .out(in_reg_wire_4[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[610]),
    .in(in_reg_wire_3[98]),
    .out(in_reg_wire_4[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[611]),
    .in(in_reg_wire_3[99]),
    .out(in_reg_wire_4[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[612]),
    .in(in_reg_wire_3[100]),
    .out(in_reg_wire_4[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[613]),
    .in(in_reg_wire_3[101]),
    .out(in_reg_wire_4[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[614]),
    .in(in_reg_wire_3[102]),
    .out(in_reg_wire_4[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[615]),
    .in(in_reg_wire_3[103]),
    .out(in_reg_wire_4[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[616]),
    .in(in_reg_wire_3[104]),
    .out(in_reg_wire_4[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[617]),
    .in(in_reg_wire_3[105]),
    .out(in_reg_wire_4[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[618]),
    .in(in_reg_wire_3[106]),
    .out(in_reg_wire_4[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[619]),
    .in(in_reg_wire_3[107]),
    .out(in_reg_wire_4[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[620]),
    .in(in_reg_wire_3[108]),
    .out(in_reg_wire_4[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[621]),
    .in(in_reg_wire_3[109]),
    .out(in_reg_wire_4[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[622]),
    .in(in_reg_wire_3[110]),
    .out(in_reg_wire_4[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[623]),
    .in(in_reg_wire_3[111]),
    .out(in_reg_wire_4[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[624]),
    .in(in_reg_wire_3[112]),
    .out(in_reg_wire_4[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[625]),
    .in(in_reg_wire_3[113]),
    .out(in_reg_wire_4[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[626]),
    .in(in_reg_wire_3[114]),
    .out(in_reg_wire_4[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[627]),
    .in(in_reg_wire_3[115]),
    .out(in_reg_wire_4[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[628]),
    .in(in_reg_wire_3[116]),
    .out(in_reg_wire_4[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[629]),
    .in(in_reg_wire_3[117]),
    .out(in_reg_wire_4[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[630]),
    .in(in_reg_wire_3[118]),
    .out(in_reg_wire_4[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[631]),
    .in(in_reg_wire_3[119]),
    .out(in_reg_wire_4[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[632]),
    .in(in_reg_wire_3[120]),
    .out(in_reg_wire_4[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[633]),
    .in(in_reg_wire_3[121]),
    .out(in_reg_wire_4[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[634]),
    .in(in_reg_wire_3[122]),
    .out(in_reg_wire_4[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[635]),
    .in(in_reg_wire_3[123]),
    .out(in_reg_wire_4[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[636]),
    .in(in_reg_wire_3[124]),
    .out(in_reg_wire_4[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[637]),
    .in(in_reg_wire_3[125]),
    .out(in_reg_wire_4[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[638]),
    .in(in_reg_wire_3[126]),
    .out(in_reg_wire_4[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[639]),
    .in(in_reg_wire_3[127]),
    .out(in_reg_wire_4[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[640]),
    .in(in_reg_wire_3[128]),
    .out(in_reg_wire_4[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[641]),
    .in(in_reg_wire_3[129]),
    .out(in_reg_wire_4[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[642]),
    .in(in_reg_wire_3[130]),
    .out(in_reg_wire_4[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[643]),
    .in(in_reg_wire_3[131]),
    .out(in_reg_wire_4[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[644]),
    .in(in_reg_wire_3[132]),
    .out(in_reg_wire_4[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[645]),
    .in(in_reg_wire_3[133]),
    .out(in_reg_wire_4[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[646]),
    .in(in_reg_wire_3[134]),
    .out(in_reg_wire_4[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[647]),
    .in(in_reg_wire_3[135]),
    .out(in_reg_wire_4[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[648]),
    .in(in_reg_wire_3[136]),
    .out(in_reg_wire_4[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[649]),
    .in(in_reg_wire_3[137]),
    .out(in_reg_wire_4[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[650]),
    .in(in_reg_wire_3[138]),
    .out(in_reg_wire_4[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[651]),
    .in(in_reg_wire_3[139]),
    .out(in_reg_wire_4[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[652]),
    .in(in_reg_wire_3[140]),
    .out(in_reg_wire_4[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[653]),
    .in(in_reg_wire_3[141]),
    .out(in_reg_wire_4[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[654]),
    .in(in_reg_wire_3[142]),
    .out(in_reg_wire_4[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[655]),
    .in(in_reg_wire_3[143]),
    .out(in_reg_wire_4[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[656]),
    .in(in_reg_wire_3[144]),
    .out(in_reg_wire_4[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[657]),
    .in(in_reg_wire_3[145]),
    .out(in_reg_wire_4[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[658]),
    .in(in_reg_wire_3[146]),
    .out(in_reg_wire_4[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[659]),
    .in(in_reg_wire_3[147]),
    .out(in_reg_wire_4[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[660]),
    .in(in_reg_wire_3[148]),
    .out(in_reg_wire_4[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[661]),
    .in(in_reg_wire_3[149]),
    .out(in_reg_wire_4[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[662]),
    .in(in_reg_wire_3[150]),
    .out(in_reg_wire_4[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[663]),
    .in(in_reg_wire_3[151]),
    .out(in_reg_wire_4[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[664]),
    .in(in_reg_wire_3[152]),
    .out(in_reg_wire_4[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[665]),
    .in(in_reg_wire_3[153]),
    .out(in_reg_wire_4[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[666]),
    .in(in_reg_wire_3[154]),
    .out(in_reg_wire_4[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[667]),
    .in(in_reg_wire_3[155]),
    .out(in_reg_wire_4[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[668]),
    .in(in_reg_wire_3[156]),
    .out(in_reg_wire_4[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[669]),
    .in(in_reg_wire_3[157]),
    .out(in_reg_wire_4[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[670]),
    .in(in_reg_wire_3[158]),
    .out(in_reg_wire_4[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[671]),
    .in(in_reg_wire_3[159]),
    .out(in_reg_wire_4[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[672]),
    .in(in_reg_wire_3[160]),
    .out(in_reg_wire_4[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[673]),
    .in(in_reg_wire_3[161]),
    .out(in_reg_wire_4[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[674]),
    .in(in_reg_wire_3[162]),
    .out(in_reg_wire_4[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[675]),
    .in(in_reg_wire_3[163]),
    .out(in_reg_wire_4[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[676]),
    .in(in_reg_wire_3[164]),
    .out(in_reg_wire_4[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[677]),
    .in(in_reg_wire_3[165]),
    .out(in_reg_wire_4[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[678]),
    .in(in_reg_wire_3[166]),
    .out(in_reg_wire_4[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[679]),
    .in(in_reg_wire_3[167]),
    .out(in_reg_wire_4[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[680]),
    .in(in_reg_wire_3[168]),
    .out(in_reg_wire_4[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[681]),
    .in(in_reg_wire_3[169]),
    .out(in_reg_wire_4[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[682]),
    .in(in_reg_wire_3[170]),
    .out(in_reg_wire_4[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[683]),
    .in(in_reg_wire_3[171]),
    .out(in_reg_wire_4[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[684]),
    .in(in_reg_wire_3[172]),
    .out(in_reg_wire_4[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[685]),
    .in(in_reg_wire_3[173]),
    .out(in_reg_wire_4[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[686]),
    .in(in_reg_wire_3[174]),
    .out(in_reg_wire_4[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[687]),
    .in(in_reg_wire_3[175]),
    .out(in_reg_wire_4[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[688]),
    .in(in_reg_wire_3[176]),
    .out(in_reg_wire_4[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[689]),
    .in(in_reg_wire_3[177]),
    .out(in_reg_wire_4[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[690]),
    .in(in_reg_wire_3[178]),
    .out(in_reg_wire_4[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[691]),
    .in(in_reg_wire_3[179]),
    .out(in_reg_wire_4[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[692]),
    .in(in_reg_wire_3[180]),
    .out(in_reg_wire_4[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[693]),
    .in(in_reg_wire_3[181]),
    .out(in_reg_wire_4[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[694]),
    .in(in_reg_wire_3[182]),
    .out(in_reg_wire_4[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[695]),
    .in(in_reg_wire_3[183]),
    .out(in_reg_wire_4[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[696]),
    .in(in_reg_wire_3[184]),
    .out(in_reg_wire_4[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[697]),
    .in(in_reg_wire_3[185]),
    .out(in_reg_wire_4[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[698]),
    .in(in_reg_wire_3[186]),
    .out(in_reg_wire_4[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[699]),
    .in(in_reg_wire_3[187]),
    .out(in_reg_wire_4[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[700]),
    .in(in_reg_wire_3[188]),
    .out(in_reg_wire_4[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[701]),
    .in(in_reg_wire_3[189]),
    .out(in_reg_wire_4[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[702]),
    .in(in_reg_wire_3[190]),
    .out(in_reg_wire_4[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[703]),
    .in(in_reg_wire_3[191]),
    .out(in_reg_wire_4[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[704]),
    .in(in_reg_wire_3[192]),
    .out(in_reg_wire_4[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[705]),
    .in(in_reg_wire_3[193]),
    .out(in_reg_wire_4[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[706]),
    .in(in_reg_wire_3[194]),
    .out(in_reg_wire_4[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[707]),
    .in(in_reg_wire_3[195]),
    .out(in_reg_wire_4[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[708]),
    .in(in_reg_wire_3[196]),
    .out(in_reg_wire_4[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[709]),
    .in(in_reg_wire_3[197]),
    .out(in_reg_wire_4[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[710]),
    .in(in_reg_wire_3[198]),
    .out(in_reg_wire_4[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[711]),
    .in(in_reg_wire_3[199]),
    .out(in_reg_wire_4[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[712]),
    .in(in_reg_wire_3[200]),
    .out(in_reg_wire_4[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[713]),
    .in(in_reg_wire_3[201]),
    .out(in_reg_wire_4[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[714]),
    .in(in_reg_wire_3[202]),
    .out(in_reg_wire_4[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[715]),
    .in(in_reg_wire_3[203]),
    .out(in_reg_wire_4[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[716]),
    .in(in_reg_wire_3[204]),
    .out(in_reg_wire_4[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[717]),
    .in(in_reg_wire_3[205]),
    .out(in_reg_wire_4[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[718]),
    .in(in_reg_wire_3[206]),
    .out(in_reg_wire_4[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[719]),
    .in(in_reg_wire_3[207]),
    .out(in_reg_wire_4[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[720]),
    .in(in_reg_wire_3[208]),
    .out(in_reg_wire_4[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[721]),
    .in(in_reg_wire_3[209]),
    .out(in_reg_wire_4[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[722]),
    .in(in_reg_wire_3[210]),
    .out(in_reg_wire_4[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[723]),
    .in(in_reg_wire_3[211]),
    .out(in_reg_wire_4[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[724]),
    .in(in_reg_wire_3[212]),
    .out(in_reg_wire_4[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[725]),
    .in(in_reg_wire_3[213]),
    .out(in_reg_wire_4[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[726]),
    .in(in_reg_wire_3[214]),
    .out(in_reg_wire_4[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[727]),
    .in(in_reg_wire_3[215]),
    .out(in_reg_wire_4[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[728]),
    .in(in_reg_wire_3[216]),
    .out(in_reg_wire_4[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[729]),
    .in(in_reg_wire_3[217]),
    .out(in_reg_wire_4[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[730]),
    .in(in_reg_wire_3[218]),
    .out(in_reg_wire_4[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[731]),
    .in(in_reg_wire_3[219]),
    .out(in_reg_wire_4[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[732]),
    .in(in_reg_wire_3[220]),
    .out(in_reg_wire_4[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[733]),
    .in(in_reg_wire_3[221]),
    .out(in_reg_wire_4[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[734]),
    .in(in_reg_wire_3[222]),
    .out(in_reg_wire_4[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[735]),
    .in(in_reg_wire_3[223]),
    .out(in_reg_wire_4[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[736]),
    .in(in_reg_wire_3[224]),
    .out(in_reg_wire_4[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[737]),
    .in(in_reg_wire_3[225]),
    .out(in_reg_wire_4[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[738]),
    .in(in_reg_wire_3[226]),
    .out(in_reg_wire_4[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[739]),
    .in(in_reg_wire_3[227]),
    .out(in_reg_wire_4[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[740]),
    .in(in_reg_wire_3[228]),
    .out(in_reg_wire_4[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[741]),
    .in(in_reg_wire_3[229]),
    .out(in_reg_wire_4[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[742]),
    .in(in_reg_wire_3[230]),
    .out(in_reg_wire_4[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[743]),
    .in(in_reg_wire_3[231]),
    .out(in_reg_wire_4[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[744]),
    .in(in_reg_wire_3[232]),
    .out(in_reg_wire_4[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[745]),
    .in(in_reg_wire_3[233]),
    .out(in_reg_wire_4[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[746]),
    .in(in_reg_wire_3[234]),
    .out(in_reg_wire_4[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[747]),
    .in(in_reg_wire_3[235]),
    .out(in_reg_wire_4[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[748]),
    .in(in_reg_wire_3[236]),
    .out(in_reg_wire_4[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[749]),
    .in(in_reg_wire_3[237]),
    .out(in_reg_wire_4[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[750]),
    .in(in_reg_wire_3[238]),
    .out(in_reg_wire_4[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[751]),
    .in(in_reg_wire_3[239]),
    .out(in_reg_wire_4[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[752]),
    .in(in_reg_wire_3[240]),
    .out(in_reg_wire_4[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[753]),
    .in(in_reg_wire_3[241]),
    .out(in_reg_wire_4[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[754]),
    .in(in_reg_wire_3[242]),
    .out(in_reg_wire_4[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[755]),
    .in(in_reg_wire_3[243]),
    .out(in_reg_wire_4[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[756]),
    .in(in_reg_wire_3[244]),
    .out(in_reg_wire_4[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[757]),
    .in(in_reg_wire_3[245]),
    .out(in_reg_wire_4[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[758]),
    .in(in_reg_wire_3[246]),
    .out(in_reg_wire_4[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[759]),
    .in(in_reg_wire_3[247]),
    .out(in_reg_wire_4[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[760]),
    .in(in_reg_wire_3[248]),
    .out(in_reg_wire_4[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[761]),
    .in(in_reg_wire_3[249]),
    .out(in_reg_wire_4[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[762]),
    .in(in_reg_wire_3[250]),
    .out(in_reg_wire_4[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[763]),
    .in(in_reg_wire_3[251]),
    .out(in_reg_wire_4[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[764]),
    .in(in_reg_wire_3[252]),
    .out(in_reg_wire_4[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[765]),
    .in(in_reg_wire_3[253]),
    .out(in_reg_wire_4[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[766]),
    .in(in_reg_wire_3[254]),
    .out(in_reg_wire_4[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[767]),
    .in(in_reg_wire_3[255]),
    .out(in_reg_wire_4[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[768]),
    .in(in_reg_wire_5[0]),
    .out(in_reg_wire_6[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[769]),
    .in(in_reg_wire_5[1]),
    .out(in_reg_wire_6[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[770]),
    .in(in_reg_wire_5[2]),
    .out(in_reg_wire_6[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[771]),
    .in(in_reg_wire_5[3]),
    .out(in_reg_wire_6[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[772]),
    .in(in_reg_wire_5[4]),
    .out(in_reg_wire_6[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[773]),
    .in(in_reg_wire_5[5]),
    .out(in_reg_wire_6[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[774]),
    .in(in_reg_wire_5[6]),
    .out(in_reg_wire_6[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[775]),
    .in(in_reg_wire_5[7]),
    .out(in_reg_wire_6[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[776]),
    .in(in_reg_wire_5[8]),
    .out(in_reg_wire_6[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[777]),
    .in(in_reg_wire_5[9]),
    .out(in_reg_wire_6[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[778]),
    .in(in_reg_wire_5[10]),
    .out(in_reg_wire_6[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[779]),
    .in(in_reg_wire_5[11]),
    .out(in_reg_wire_6[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[780]),
    .in(in_reg_wire_5[12]),
    .out(in_reg_wire_6[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[781]),
    .in(in_reg_wire_5[13]),
    .out(in_reg_wire_6[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[782]),
    .in(in_reg_wire_5[14]),
    .out(in_reg_wire_6[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[783]),
    .in(in_reg_wire_5[15]),
    .out(in_reg_wire_6[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[784]),
    .in(in_reg_wire_5[16]),
    .out(in_reg_wire_6[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[785]),
    .in(in_reg_wire_5[17]),
    .out(in_reg_wire_6[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[786]),
    .in(in_reg_wire_5[18]),
    .out(in_reg_wire_6[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[787]),
    .in(in_reg_wire_5[19]),
    .out(in_reg_wire_6[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[788]),
    .in(in_reg_wire_5[20]),
    .out(in_reg_wire_6[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[789]),
    .in(in_reg_wire_5[21]),
    .out(in_reg_wire_6[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[790]),
    .in(in_reg_wire_5[22]),
    .out(in_reg_wire_6[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[791]),
    .in(in_reg_wire_5[23]),
    .out(in_reg_wire_6[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[792]),
    .in(in_reg_wire_5[24]),
    .out(in_reg_wire_6[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[793]),
    .in(in_reg_wire_5[25]),
    .out(in_reg_wire_6[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[794]),
    .in(in_reg_wire_5[26]),
    .out(in_reg_wire_6[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[795]),
    .in(in_reg_wire_5[27]),
    .out(in_reg_wire_6[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[796]),
    .in(in_reg_wire_5[28]),
    .out(in_reg_wire_6[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[797]),
    .in(in_reg_wire_5[29]),
    .out(in_reg_wire_6[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[798]),
    .in(in_reg_wire_5[30]),
    .out(in_reg_wire_6[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[799]),
    .in(in_reg_wire_5[31]),
    .out(in_reg_wire_6[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[800]),
    .in(in_reg_wire_5[32]),
    .out(in_reg_wire_6[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[801]),
    .in(in_reg_wire_5[33]),
    .out(in_reg_wire_6[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[802]),
    .in(in_reg_wire_5[34]),
    .out(in_reg_wire_6[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[803]),
    .in(in_reg_wire_5[35]),
    .out(in_reg_wire_6[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[804]),
    .in(in_reg_wire_5[36]),
    .out(in_reg_wire_6[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[805]),
    .in(in_reg_wire_5[37]),
    .out(in_reg_wire_6[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[806]),
    .in(in_reg_wire_5[38]),
    .out(in_reg_wire_6[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[807]),
    .in(in_reg_wire_5[39]),
    .out(in_reg_wire_6[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[808]),
    .in(in_reg_wire_5[40]),
    .out(in_reg_wire_6[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[809]),
    .in(in_reg_wire_5[41]),
    .out(in_reg_wire_6[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[810]),
    .in(in_reg_wire_5[42]),
    .out(in_reg_wire_6[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[811]),
    .in(in_reg_wire_5[43]),
    .out(in_reg_wire_6[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[812]),
    .in(in_reg_wire_5[44]),
    .out(in_reg_wire_6[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[813]),
    .in(in_reg_wire_5[45]),
    .out(in_reg_wire_6[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[814]),
    .in(in_reg_wire_5[46]),
    .out(in_reg_wire_6[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[815]),
    .in(in_reg_wire_5[47]),
    .out(in_reg_wire_6[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[816]),
    .in(in_reg_wire_5[48]),
    .out(in_reg_wire_6[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[817]),
    .in(in_reg_wire_5[49]),
    .out(in_reg_wire_6[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[818]),
    .in(in_reg_wire_5[50]),
    .out(in_reg_wire_6[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[819]),
    .in(in_reg_wire_5[51]),
    .out(in_reg_wire_6[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[820]),
    .in(in_reg_wire_5[52]),
    .out(in_reg_wire_6[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[821]),
    .in(in_reg_wire_5[53]),
    .out(in_reg_wire_6[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[822]),
    .in(in_reg_wire_5[54]),
    .out(in_reg_wire_6[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[823]),
    .in(in_reg_wire_5[55]),
    .out(in_reg_wire_6[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[824]),
    .in(in_reg_wire_5[56]),
    .out(in_reg_wire_6[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[825]),
    .in(in_reg_wire_5[57]),
    .out(in_reg_wire_6[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[826]),
    .in(in_reg_wire_5[58]),
    .out(in_reg_wire_6[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[827]),
    .in(in_reg_wire_5[59]),
    .out(in_reg_wire_6[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[828]),
    .in(in_reg_wire_5[60]),
    .out(in_reg_wire_6[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[829]),
    .in(in_reg_wire_5[61]),
    .out(in_reg_wire_6[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[830]),
    .in(in_reg_wire_5[62]),
    .out(in_reg_wire_6[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[831]),
    .in(in_reg_wire_5[63]),
    .out(in_reg_wire_6[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[832]),
    .in(in_reg_wire_5[64]),
    .out(in_reg_wire_6[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[833]),
    .in(in_reg_wire_5[65]),
    .out(in_reg_wire_6[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[834]),
    .in(in_reg_wire_5[66]),
    .out(in_reg_wire_6[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[835]),
    .in(in_reg_wire_5[67]),
    .out(in_reg_wire_6[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[836]),
    .in(in_reg_wire_5[68]),
    .out(in_reg_wire_6[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[837]),
    .in(in_reg_wire_5[69]),
    .out(in_reg_wire_6[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[838]),
    .in(in_reg_wire_5[70]),
    .out(in_reg_wire_6[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[839]),
    .in(in_reg_wire_5[71]),
    .out(in_reg_wire_6[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[840]),
    .in(in_reg_wire_5[72]),
    .out(in_reg_wire_6[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[841]),
    .in(in_reg_wire_5[73]),
    .out(in_reg_wire_6[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[842]),
    .in(in_reg_wire_5[74]),
    .out(in_reg_wire_6[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[843]),
    .in(in_reg_wire_5[75]),
    .out(in_reg_wire_6[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[844]),
    .in(in_reg_wire_5[76]),
    .out(in_reg_wire_6[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[845]),
    .in(in_reg_wire_5[77]),
    .out(in_reg_wire_6[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[846]),
    .in(in_reg_wire_5[78]),
    .out(in_reg_wire_6[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[847]),
    .in(in_reg_wire_5[79]),
    .out(in_reg_wire_6[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[848]),
    .in(in_reg_wire_5[80]),
    .out(in_reg_wire_6[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[849]),
    .in(in_reg_wire_5[81]),
    .out(in_reg_wire_6[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[850]),
    .in(in_reg_wire_5[82]),
    .out(in_reg_wire_6[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[851]),
    .in(in_reg_wire_5[83]),
    .out(in_reg_wire_6[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[852]),
    .in(in_reg_wire_5[84]),
    .out(in_reg_wire_6[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[853]),
    .in(in_reg_wire_5[85]),
    .out(in_reg_wire_6[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[854]),
    .in(in_reg_wire_5[86]),
    .out(in_reg_wire_6[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[855]),
    .in(in_reg_wire_5[87]),
    .out(in_reg_wire_6[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[856]),
    .in(in_reg_wire_5[88]),
    .out(in_reg_wire_6[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[857]),
    .in(in_reg_wire_5[89]),
    .out(in_reg_wire_6[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[858]),
    .in(in_reg_wire_5[90]),
    .out(in_reg_wire_6[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[859]),
    .in(in_reg_wire_5[91]),
    .out(in_reg_wire_6[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[860]),
    .in(in_reg_wire_5[92]),
    .out(in_reg_wire_6[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[861]),
    .in(in_reg_wire_5[93]),
    .out(in_reg_wire_6[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[862]),
    .in(in_reg_wire_5[94]),
    .out(in_reg_wire_6[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[863]),
    .in(in_reg_wire_5[95]),
    .out(in_reg_wire_6[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[864]),
    .in(in_reg_wire_5[96]),
    .out(in_reg_wire_6[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[865]),
    .in(in_reg_wire_5[97]),
    .out(in_reg_wire_6[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[866]),
    .in(in_reg_wire_5[98]),
    .out(in_reg_wire_6[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[867]),
    .in(in_reg_wire_5[99]),
    .out(in_reg_wire_6[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[868]),
    .in(in_reg_wire_5[100]),
    .out(in_reg_wire_6[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[869]),
    .in(in_reg_wire_5[101]),
    .out(in_reg_wire_6[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[870]),
    .in(in_reg_wire_5[102]),
    .out(in_reg_wire_6[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[871]),
    .in(in_reg_wire_5[103]),
    .out(in_reg_wire_6[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[872]),
    .in(in_reg_wire_5[104]),
    .out(in_reg_wire_6[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[873]),
    .in(in_reg_wire_5[105]),
    .out(in_reg_wire_6[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[874]),
    .in(in_reg_wire_5[106]),
    .out(in_reg_wire_6[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[875]),
    .in(in_reg_wire_5[107]),
    .out(in_reg_wire_6[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[876]),
    .in(in_reg_wire_5[108]),
    .out(in_reg_wire_6[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[877]),
    .in(in_reg_wire_5[109]),
    .out(in_reg_wire_6[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[878]),
    .in(in_reg_wire_5[110]),
    .out(in_reg_wire_6[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[879]),
    .in(in_reg_wire_5[111]),
    .out(in_reg_wire_6[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[880]),
    .in(in_reg_wire_5[112]),
    .out(in_reg_wire_6[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[881]),
    .in(in_reg_wire_5[113]),
    .out(in_reg_wire_6[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[882]),
    .in(in_reg_wire_5[114]),
    .out(in_reg_wire_6[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[883]),
    .in(in_reg_wire_5[115]),
    .out(in_reg_wire_6[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[884]),
    .in(in_reg_wire_5[116]),
    .out(in_reg_wire_6[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[885]),
    .in(in_reg_wire_5[117]),
    .out(in_reg_wire_6[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[886]),
    .in(in_reg_wire_5[118]),
    .out(in_reg_wire_6[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[887]),
    .in(in_reg_wire_5[119]),
    .out(in_reg_wire_6[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[888]),
    .in(in_reg_wire_5[120]),
    .out(in_reg_wire_6[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[889]),
    .in(in_reg_wire_5[121]),
    .out(in_reg_wire_6[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[890]),
    .in(in_reg_wire_5[122]),
    .out(in_reg_wire_6[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[891]),
    .in(in_reg_wire_5[123]),
    .out(in_reg_wire_6[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[892]),
    .in(in_reg_wire_5[124]),
    .out(in_reg_wire_6[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[893]),
    .in(in_reg_wire_5[125]),
    .out(in_reg_wire_6[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[894]),
    .in(in_reg_wire_5[126]),
    .out(in_reg_wire_6[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[895]),
    .in(in_reg_wire_5[127]),
    .out(in_reg_wire_6[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[896]),
    .in(in_reg_wire_5[128]),
    .out(in_reg_wire_6[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[897]),
    .in(in_reg_wire_5[129]),
    .out(in_reg_wire_6[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[898]),
    .in(in_reg_wire_5[130]),
    .out(in_reg_wire_6[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[899]),
    .in(in_reg_wire_5[131]),
    .out(in_reg_wire_6[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[900]),
    .in(in_reg_wire_5[132]),
    .out(in_reg_wire_6[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[901]),
    .in(in_reg_wire_5[133]),
    .out(in_reg_wire_6[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[902]),
    .in(in_reg_wire_5[134]),
    .out(in_reg_wire_6[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[903]),
    .in(in_reg_wire_5[135]),
    .out(in_reg_wire_6[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[904]),
    .in(in_reg_wire_5[136]),
    .out(in_reg_wire_6[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[905]),
    .in(in_reg_wire_5[137]),
    .out(in_reg_wire_6[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[906]),
    .in(in_reg_wire_5[138]),
    .out(in_reg_wire_6[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[907]),
    .in(in_reg_wire_5[139]),
    .out(in_reg_wire_6[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[908]),
    .in(in_reg_wire_5[140]),
    .out(in_reg_wire_6[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[909]),
    .in(in_reg_wire_5[141]),
    .out(in_reg_wire_6[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[910]),
    .in(in_reg_wire_5[142]),
    .out(in_reg_wire_6[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[911]),
    .in(in_reg_wire_5[143]),
    .out(in_reg_wire_6[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[912]),
    .in(in_reg_wire_5[144]),
    .out(in_reg_wire_6[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[913]),
    .in(in_reg_wire_5[145]),
    .out(in_reg_wire_6[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[914]),
    .in(in_reg_wire_5[146]),
    .out(in_reg_wire_6[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[915]),
    .in(in_reg_wire_5[147]),
    .out(in_reg_wire_6[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[916]),
    .in(in_reg_wire_5[148]),
    .out(in_reg_wire_6[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[917]),
    .in(in_reg_wire_5[149]),
    .out(in_reg_wire_6[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[918]),
    .in(in_reg_wire_5[150]),
    .out(in_reg_wire_6[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[919]),
    .in(in_reg_wire_5[151]),
    .out(in_reg_wire_6[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[920]),
    .in(in_reg_wire_5[152]),
    .out(in_reg_wire_6[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[921]),
    .in(in_reg_wire_5[153]),
    .out(in_reg_wire_6[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[922]),
    .in(in_reg_wire_5[154]),
    .out(in_reg_wire_6[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[923]),
    .in(in_reg_wire_5[155]),
    .out(in_reg_wire_6[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[924]),
    .in(in_reg_wire_5[156]),
    .out(in_reg_wire_6[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[925]),
    .in(in_reg_wire_5[157]),
    .out(in_reg_wire_6[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[926]),
    .in(in_reg_wire_5[158]),
    .out(in_reg_wire_6[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[927]),
    .in(in_reg_wire_5[159]),
    .out(in_reg_wire_6[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[928]),
    .in(in_reg_wire_5[160]),
    .out(in_reg_wire_6[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[929]),
    .in(in_reg_wire_5[161]),
    .out(in_reg_wire_6[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[930]),
    .in(in_reg_wire_5[162]),
    .out(in_reg_wire_6[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[931]),
    .in(in_reg_wire_5[163]),
    .out(in_reg_wire_6[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[932]),
    .in(in_reg_wire_5[164]),
    .out(in_reg_wire_6[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[933]),
    .in(in_reg_wire_5[165]),
    .out(in_reg_wire_6[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[934]),
    .in(in_reg_wire_5[166]),
    .out(in_reg_wire_6[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[935]),
    .in(in_reg_wire_5[167]),
    .out(in_reg_wire_6[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[936]),
    .in(in_reg_wire_5[168]),
    .out(in_reg_wire_6[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[937]),
    .in(in_reg_wire_5[169]),
    .out(in_reg_wire_6[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[938]),
    .in(in_reg_wire_5[170]),
    .out(in_reg_wire_6[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[939]),
    .in(in_reg_wire_5[171]),
    .out(in_reg_wire_6[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[940]),
    .in(in_reg_wire_5[172]),
    .out(in_reg_wire_6[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[941]),
    .in(in_reg_wire_5[173]),
    .out(in_reg_wire_6[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[942]),
    .in(in_reg_wire_5[174]),
    .out(in_reg_wire_6[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[943]),
    .in(in_reg_wire_5[175]),
    .out(in_reg_wire_6[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[944]),
    .in(in_reg_wire_5[176]),
    .out(in_reg_wire_6[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[945]),
    .in(in_reg_wire_5[177]),
    .out(in_reg_wire_6[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[946]),
    .in(in_reg_wire_5[178]),
    .out(in_reg_wire_6[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[947]),
    .in(in_reg_wire_5[179]),
    .out(in_reg_wire_6[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[948]),
    .in(in_reg_wire_5[180]),
    .out(in_reg_wire_6[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[949]),
    .in(in_reg_wire_5[181]),
    .out(in_reg_wire_6[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[950]),
    .in(in_reg_wire_5[182]),
    .out(in_reg_wire_6[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[951]),
    .in(in_reg_wire_5[183]),
    .out(in_reg_wire_6[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[952]),
    .in(in_reg_wire_5[184]),
    .out(in_reg_wire_6[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[953]),
    .in(in_reg_wire_5[185]),
    .out(in_reg_wire_6[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[954]),
    .in(in_reg_wire_5[186]),
    .out(in_reg_wire_6[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[955]),
    .in(in_reg_wire_5[187]),
    .out(in_reg_wire_6[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[956]),
    .in(in_reg_wire_5[188]),
    .out(in_reg_wire_6[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[957]),
    .in(in_reg_wire_5[189]),
    .out(in_reg_wire_6[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[958]),
    .in(in_reg_wire_5[190]),
    .out(in_reg_wire_6[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[959]),
    .in(in_reg_wire_5[191]),
    .out(in_reg_wire_6[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[960]),
    .in(in_reg_wire_5[192]),
    .out(in_reg_wire_6[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[961]),
    .in(in_reg_wire_5[193]),
    .out(in_reg_wire_6[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[962]),
    .in(in_reg_wire_5[194]),
    .out(in_reg_wire_6[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[963]),
    .in(in_reg_wire_5[195]),
    .out(in_reg_wire_6[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[964]),
    .in(in_reg_wire_5[196]),
    .out(in_reg_wire_6[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[965]),
    .in(in_reg_wire_5[197]),
    .out(in_reg_wire_6[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[966]),
    .in(in_reg_wire_5[198]),
    .out(in_reg_wire_6[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[967]),
    .in(in_reg_wire_5[199]),
    .out(in_reg_wire_6[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[968]),
    .in(in_reg_wire_5[200]),
    .out(in_reg_wire_6[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[969]),
    .in(in_reg_wire_5[201]),
    .out(in_reg_wire_6[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[970]),
    .in(in_reg_wire_5[202]),
    .out(in_reg_wire_6[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[971]),
    .in(in_reg_wire_5[203]),
    .out(in_reg_wire_6[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[972]),
    .in(in_reg_wire_5[204]),
    .out(in_reg_wire_6[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[973]),
    .in(in_reg_wire_5[205]),
    .out(in_reg_wire_6[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[974]),
    .in(in_reg_wire_5[206]),
    .out(in_reg_wire_6[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[975]),
    .in(in_reg_wire_5[207]),
    .out(in_reg_wire_6[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[976]),
    .in(in_reg_wire_5[208]),
    .out(in_reg_wire_6[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[977]),
    .in(in_reg_wire_5[209]),
    .out(in_reg_wire_6[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[978]),
    .in(in_reg_wire_5[210]),
    .out(in_reg_wire_6[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[979]),
    .in(in_reg_wire_5[211]),
    .out(in_reg_wire_6[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[980]),
    .in(in_reg_wire_5[212]),
    .out(in_reg_wire_6[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[981]),
    .in(in_reg_wire_5[213]),
    .out(in_reg_wire_6[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[982]),
    .in(in_reg_wire_5[214]),
    .out(in_reg_wire_6[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[983]),
    .in(in_reg_wire_5[215]),
    .out(in_reg_wire_6[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[984]),
    .in(in_reg_wire_5[216]),
    .out(in_reg_wire_6[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[985]),
    .in(in_reg_wire_5[217]),
    .out(in_reg_wire_6[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[986]),
    .in(in_reg_wire_5[218]),
    .out(in_reg_wire_6[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[987]),
    .in(in_reg_wire_5[219]),
    .out(in_reg_wire_6[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[988]),
    .in(in_reg_wire_5[220]),
    .out(in_reg_wire_6[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[989]),
    .in(in_reg_wire_5[221]),
    .out(in_reg_wire_6[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[990]),
    .in(in_reg_wire_5[222]),
    .out(in_reg_wire_6[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[991]),
    .in(in_reg_wire_5[223]),
    .out(in_reg_wire_6[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[992]),
    .in(in_reg_wire_5[224]),
    .out(in_reg_wire_6[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[993]),
    .in(in_reg_wire_5[225]),
    .out(in_reg_wire_6[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[994]),
    .in(in_reg_wire_5[226]),
    .out(in_reg_wire_6[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[995]),
    .in(in_reg_wire_5[227]),
    .out(in_reg_wire_6[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[996]),
    .in(in_reg_wire_5[228]),
    .out(in_reg_wire_6[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[997]),
    .in(in_reg_wire_5[229]),
    .out(in_reg_wire_6[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[998]),
    .in(in_reg_wire_5[230]),
    .out(in_reg_wire_6[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[999]),
    .in(in_reg_wire_5[231]),
    .out(in_reg_wire_6[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1000]),
    .in(in_reg_wire_5[232]),
    .out(in_reg_wire_6[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1001]),
    .in(in_reg_wire_5[233]),
    .out(in_reg_wire_6[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1002]),
    .in(in_reg_wire_5[234]),
    .out(in_reg_wire_6[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1003]),
    .in(in_reg_wire_5[235]),
    .out(in_reg_wire_6[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1004]),
    .in(in_reg_wire_5[236]),
    .out(in_reg_wire_6[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1005]),
    .in(in_reg_wire_5[237]),
    .out(in_reg_wire_6[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1006]),
    .in(in_reg_wire_5[238]),
    .out(in_reg_wire_6[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1007]),
    .in(in_reg_wire_5[239]),
    .out(in_reg_wire_6[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1008]),
    .in(in_reg_wire_5[240]),
    .out(in_reg_wire_6[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1009]),
    .in(in_reg_wire_5[241]),
    .out(in_reg_wire_6[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1010]),
    .in(in_reg_wire_5[242]),
    .out(in_reg_wire_6[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1011]),
    .in(in_reg_wire_5[243]),
    .out(in_reg_wire_6[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1012]),
    .in(in_reg_wire_5[244]),
    .out(in_reg_wire_6[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1013]),
    .in(in_reg_wire_5[245]),
    .out(in_reg_wire_6[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1014]),
    .in(in_reg_wire_5[246]),
    .out(in_reg_wire_6[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1015]),
    .in(in_reg_wire_5[247]),
    .out(in_reg_wire_6[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1016]),
    .in(in_reg_wire_5[248]),
    .out(in_reg_wire_6[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1017]),
    .in(in_reg_wire_5[249]),
    .out(in_reg_wire_6[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1018]),
    .in(in_reg_wire_5[250]),
    .out(in_reg_wire_6[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1019]),
    .in(in_reg_wire_5[251]),
    .out(in_reg_wire_6[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1020]),
    .in(in_reg_wire_5[252]),
    .out(in_reg_wire_6[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1021]),
    .in(in_reg_wire_5[253]),
    .out(in_reg_wire_6[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1022]),
    .in(in_reg_wire_5[254]),
    .out(in_reg_wire_6[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1023]),
    .in(in_reg_wire_5[255]),
    .out(in_reg_wire_6[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1024]),
    .in(in_reg_wire_7[0]),
    .out(out0)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1025]),
    .in(in_reg_wire_7[1]),
    .out(out4)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1026]),
    .in(in_reg_wire_7[2]),
    .out(out8)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1027]),
    .in(in_reg_wire_7[3]),
    .out(out12)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1028]),
    .in(in_reg_wire_7[4]),
    .out(out16)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1029]),
    .in(in_reg_wire_7[5]),
    .out(out20)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1030]),
    .in(in_reg_wire_7[6]),
    .out(out24)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1031]),
    .in(in_reg_wire_7[7]),
    .out(out28)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1032]),
    .in(in_reg_wire_7[8]),
    .out(out32)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1033]),
    .in(in_reg_wire_7[9]),
    .out(out36)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1034]),
    .in(in_reg_wire_7[10]),
    .out(out40)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1035]),
    .in(in_reg_wire_7[11]),
    .out(out44)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1036]),
    .in(in_reg_wire_7[12]),
    .out(out48)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1037]),
    .in(in_reg_wire_7[13]),
    .out(out52)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1038]),
    .in(in_reg_wire_7[14]),
    .out(out56)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1039]),
    .in(in_reg_wire_7[15]),
    .out(out60)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1040]),
    .in(in_reg_wire_7[16]),
    .out(out64)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1041]),
    .in(in_reg_wire_7[17]),
    .out(out68)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1042]),
    .in(in_reg_wire_7[18]),
    .out(out72)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1043]),
    .in(in_reg_wire_7[19]),
    .out(out76)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1044]),
    .in(in_reg_wire_7[20]),
    .out(out80)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1045]),
    .in(in_reg_wire_7[21]),
    .out(out84)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1046]),
    .in(in_reg_wire_7[22]),
    .out(out88)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1047]),
    .in(in_reg_wire_7[23]),
    .out(out92)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1048]),
    .in(in_reg_wire_7[24]),
    .out(out96)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1049]),
    .in(in_reg_wire_7[25]),
    .out(out100)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1050]),
    .in(in_reg_wire_7[26]),
    .out(out104)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1051]),
    .in(in_reg_wire_7[27]),
    .out(out108)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1052]),
    .in(in_reg_wire_7[28]),
    .out(out112)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1053]),
    .in(in_reg_wire_7[29]),
    .out(out116)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1054]),
    .in(in_reg_wire_7[30]),
    .out(out120)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1055]),
    .in(in_reg_wire_7[31]),
    .out(out124)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1056]),
    .in(in_reg_wire_7[32]),
    .out(out128)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1057]),
    .in(in_reg_wire_7[33]),
    .out(out132)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1058]),
    .in(in_reg_wire_7[34]),
    .out(out136)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1059]),
    .in(in_reg_wire_7[35]),
    .out(out140)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1060]),
    .in(in_reg_wire_7[36]),
    .out(out144)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1061]),
    .in(in_reg_wire_7[37]),
    .out(out148)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1062]),
    .in(in_reg_wire_7[38]),
    .out(out152)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1063]),
    .in(in_reg_wire_7[39]),
    .out(out156)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1064]),
    .in(in_reg_wire_7[40]),
    .out(out160)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1065]),
    .in(in_reg_wire_7[41]),
    .out(out164)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1066]),
    .in(in_reg_wire_7[42]),
    .out(out168)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1067]),
    .in(in_reg_wire_7[43]),
    .out(out172)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1068]),
    .in(in_reg_wire_7[44]),
    .out(out176)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1069]),
    .in(in_reg_wire_7[45]),
    .out(out180)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1070]),
    .in(in_reg_wire_7[46]),
    .out(out184)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1071]),
    .in(in_reg_wire_7[47]),
    .out(out188)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1072]),
    .in(in_reg_wire_7[48]),
    .out(out192)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1073]),
    .in(in_reg_wire_7[49]),
    .out(out196)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1074]),
    .in(in_reg_wire_7[50]),
    .out(out200)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1075]),
    .in(in_reg_wire_7[51]),
    .out(out204)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1076]),
    .in(in_reg_wire_7[52]),
    .out(out208)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1077]),
    .in(in_reg_wire_7[53]),
    .out(out212)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1078]),
    .in(in_reg_wire_7[54]),
    .out(out216)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1079]),
    .in(in_reg_wire_7[55]),
    .out(out220)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1080]),
    .in(in_reg_wire_7[56]),
    .out(out224)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1081]),
    .in(in_reg_wire_7[57]),
    .out(out228)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1082]),
    .in(in_reg_wire_7[58]),
    .out(out232)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1083]),
    .in(in_reg_wire_7[59]),
    .out(out236)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1084]),
    .in(in_reg_wire_7[60]),
    .out(out240)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1085]),
    .in(in_reg_wire_7[61]),
    .out(out244)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1086]),
    .in(in_reg_wire_7[62]),
    .out(out248)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1087]),
    .in(in_reg_wire_7[63]),
    .out(out252)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1088]),
    .in(in_reg_wire_7[64]),
    .out(out1)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1089]),
    .in(in_reg_wire_7[65]),
    .out(out5)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1090]),
    .in(in_reg_wire_7[66]),
    .out(out9)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1091]),
    .in(in_reg_wire_7[67]),
    .out(out13)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1092]),
    .in(in_reg_wire_7[68]),
    .out(out17)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1093]),
    .in(in_reg_wire_7[69]),
    .out(out21)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1094]),
    .in(in_reg_wire_7[70]),
    .out(out25)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1095]),
    .in(in_reg_wire_7[71]),
    .out(out29)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1096]),
    .in(in_reg_wire_7[72]),
    .out(out33)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1097]),
    .in(in_reg_wire_7[73]),
    .out(out37)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1098]),
    .in(in_reg_wire_7[74]),
    .out(out41)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1099]),
    .in(in_reg_wire_7[75]),
    .out(out45)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1100]),
    .in(in_reg_wire_7[76]),
    .out(out49)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1101]),
    .in(in_reg_wire_7[77]),
    .out(out53)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1102]),
    .in(in_reg_wire_7[78]),
    .out(out57)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1103]),
    .in(in_reg_wire_7[79]),
    .out(out61)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1104]),
    .in(in_reg_wire_7[80]),
    .out(out65)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1105]),
    .in(in_reg_wire_7[81]),
    .out(out69)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1106]),
    .in(in_reg_wire_7[82]),
    .out(out73)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1107]),
    .in(in_reg_wire_7[83]),
    .out(out77)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1108]),
    .in(in_reg_wire_7[84]),
    .out(out81)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1109]),
    .in(in_reg_wire_7[85]),
    .out(out85)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1110]),
    .in(in_reg_wire_7[86]),
    .out(out89)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1111]),
    .in(in_reg_wire_7[87]),
    .out(out93)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1112]),
    .in(in_reg_wire_7[88]),
    .out(out97)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1113]),
    .in(in_reg_wire_7[89]),
    .out(out101)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1114]),
    .in(in_reg_wire_7[90]),
    .out(out105)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1115]),
    .in(in_reg_wire_7[91]),
    .out(out109)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1116]),
    .in(in_reg_wire_7[92]),
    .out(out113)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1117]),
    .in(in_reg_wire_7[93]),
    .out(out117)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1118]),
    .in(in_reg_wire_7[94]),
    .out(out121)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1119]),
    .in(in_reg_wire_7[95]),
    .out(out125)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1120]),
    .in(in_reg_wire_7[96]),
    .out(out129)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1121]),
    .in(in_reg_wire_7[97]),
    .out(out133)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1122]),
    .in(in_reg_wire_7[98]),
    .out(out137)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1123]),
    .in(in_reg_wire_7[99]),
    .out(out141)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1124]),
    .in(in_reg_wire_7[100]),
    .out(out145)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1125]),
    .in(in_reg_wire_7[101]),
    .out(out149)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1126]),
    .in(in_reg_wire_7[102]),
    .out(out153)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1127]),
    .in(in_reg_wire_7[103]),
    .out(out157)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1128]),
    .in(in_reg_wire_7[104]),
    .out(out161)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1129]),
    .in(in_reg_wire_7[105]),
    .out(out165)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1130]),
    .in(in_reg_wire_7[106]),
    .out(out169)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1131]),
    .in(in_reg_wire_7[107]),
    .out(out173)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1132]),
    .in(in_reg_wire_7[108]),
    .out(out177)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1133]),
    .in(in_reg_wire_7[109]),
    .out(out181)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1134]),
    .in(in_reg_wire_7[110]),
    .out(out185)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1135]),
    .in(in_reg_wire_7[111]),
    .out(out189)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1136]),
    .in(in_reg_wire_7[112]),
    .out(out193)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1137]),
    .in(in_reg_wire_7[113]),
    .out(out197)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1138]),
    .in(in_reg_wire_7[114]),
    .out(out201)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1139]),
    .in(in_reg_wire_7[115]),
    .out(out205)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1140]),
    .in(in_reg_wire_7[116]),
    .out(out209)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1141]),
    .in(in_reg_wire_7[117]),
    .out(out213)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1142]),
    .in(in_reg_wire_7[118]),
    .out(out217)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1143]),
    .in(in_reg_wire_7[119]),
    .out(out221)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1144]),
    .in(in_reg_wire_7[120]),
    .out(out225)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1145]),
    .in(in_reg_wire_7[121]),
    .out(out229)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1146]),
    .in(in_reg_wire_7[122]),
    .out(out233)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1147]),
    .in(in_reg_wire_7[123]),
    .out(out237)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1148]),
    .in(in_reg_wire_7[124]),
    .out(out241)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1149]),
    .in(in_reg_wire_7[125]),
    .out(out245)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1150]),
    .in(in_reg_wire_7[126]),
    .out(out249)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1151]),
    .in(in_reg_wire_7[127]),
    .out(out253)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1152]),
    .in(in_reg_wire_7[128]),
    .out(out2)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1153]),
    .in(in_reg_wire_7[129]),
    .out(out6)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1154]),
    .in(in_reg_wire_7[130]),
    .out(out10)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1155]),
    .in(in_reg_wire_7[131]),
    .out(out14)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1156]),
    .in(in_reg_wire_7[132]),
    .out(out18)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1157]),
    .in(in_reg_wire_7[133]),
    .out(out22)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1158]),
    .in(in_reg_wire_7[134]),
    .out(out26)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1159]),
    .in(in_reg_wire_7[135]),
    .out(out30)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1160]),
    .in(in_reg_wire_7[136]),
    .out(out34)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1161]),
    .in(in_reg_wire_7[137]),
    .out(out38)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1162]),
    .in(in_reg_wire_7[138]),
    .out(out42)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1163]),
    .in(in_reg_wire_7[139]),
    .out(out46)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1164]),
    .in(in_reg_wire_7[140]),
    .out(out50)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1165]),
    .in(in_reg_wire_7[141]),
    .out(out54)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1166]),
    .in(in_reg_wire_7[142]),
    .out(out58)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1167]),
    .in(in_reg_wire_7[143]),
    .out(out62)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1168]),
    .in(in_reg_wire_7[144]),
    .out(out66)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1169]),
    .in(in_reg_wire_7[145]),
    .out(out70)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1170]),
    .in(in_reg_wire_7[146]),
    .out(out74)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1171]),
    .in(in_reg_wire_7[147]),
    .out(out78)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1172]),
    .in(in_reg_wire_7[148]),
    .out(out82)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1173]),
    .in(in_reg_wire_7[149]),
    .out(out86)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1174]),
    .in(in_reg_wire_7[150]),
    .out(out90)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1175]),
    .in(in_reg_wire_7[151]),
    .out(out94)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1176]),
    .in(in_reg_wire_7[152]),
    .out(out98)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1177]),
    .in(in_reg_wire_7[153]),
    .out(out102)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1178]),
    .in(in_reg_wire_7[154]),
    .out(out106)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1179]),
    .in(in_reg_wire_7[155]),
    .out(out110)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1180]),
    .in(in_reg_wire_7[156]),
    .out(out114)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1181]),
    .in(in_reg_wire_7[157]),
    .out(out118)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1182]),
    .in(in_reg_wire_7[158]),
    .out(out122)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1183]),
    .in(in_reg_wire_7[159]),
    .out(out126)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1184]),
    .in(in_reg_wire_7[160]),
    .out(out130)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1185]),
    .in(in_reg_wire_7[161]),
    .out(out134)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1186]),
    .in(in_reg_wire_7[162]),
    .out(out138)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1187]),
    .in(in_reg_wire_7[163]),
    .out(out142)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1188]),
    .in(in_reg_wire_7[164]),
    .out(out146)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1189]),
    .in(in_reg_wire_7[165]),
    .out(out150)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1190]),
    .in(in_reg_wire_7[166]),
    .out(out154)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1191]),
    .in(in_reg_wire_7[167]),
    .out(out158)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1192]),
    .in(in_reg_wire_7[168]),
    .out(out162)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1193]),
    .in(in_reg_wire_7[169]),
    .out(out166)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1194]),
    .in(in_reg_wire_7[170]),
    .out(out170)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1195]),
    .in(in_reg_wire_7[171]),
    .out(out174)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1196]),
    .in(in_reg_wire_7[172]),
    .out(out178)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1197]),
    .in(in_reg_wire_7[173]),
    .out(out182)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1198]),
    .in(in_reg_wire_7[174]),
    .out(out186)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1199]),
    .in(in_reg_wire_7[175]),
    .out(out190)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1200]),
    .in(in_reg_wire_7[176]),
    .out(out194)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1201]),
    .in(in_reg_wire_7[177]),
    .out(out198)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1202]),
    .in(in_reg_wire_7[178]),
    .out(out202)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1203]),
    .in(in_reg_wire_7[179]),
    .out(out206)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1204]),
    .in(in_reg_wire_7[180]),
    .out(out210)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1205]),
    .in(in_reg_wire_7[181]),
    .out(out214)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1206]),
    .in(in_reg_wire_7[182]),
    .out(out218)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1207]),
    .in(in_reg_wire_7[183]),
    .out(out222)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1208]),
    .in(in_reg_wire_7[184]),
    .out(out226)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1209]),
    .in(in_reg_wire_7[185]),
    .out(out230)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1210]),
    .in(in_reg_wire_7[186]),
    .out(out234)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1211]),
    .in(in_reg_wire_7[187]),
    .out(out238)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1212]),
    .in(in_reg_wire_7[188]),
    .out(out242)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1213]),
    .in(in_reg_wire_7[189]),
    .out(out246)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1214]),
    .in(in_reg_wire_7[190]),
    .out(out250)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1215]),
    .in(in_reg_wire_7[191]),
    .out(out254)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1216]),
    .in(in_reg_wire_7[192]),
    .out(out3)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1217]),
    .in(in_reg_wire_7[193]),
    .out(out7)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1218]),
    .in(in_reg_wire_7[194]),
    .out(out11)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1219]),
    .in(in_reg_wire_7[195]),
    .out(out15)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1220]),
    .in(in_reg_wire_7[196]),
    .out(out19)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1221]),
    .in(in_reg_wire_7[197]),
    .out(out23)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1222]),
    .in(in_reg_wire_7[198]),
    .out(out27)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1223]),
    .in(in_reg_wire_7[199]),
    .out(out31)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1224]),
    .in(in_reg_wire_7[200]),
    .out(out35)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1225]),
    .in(in_reg_wire_7[201]),
    .out(out39)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1226]),
    .in(in_reg_wire_7[202]),
    .out(out43)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1227]),
    .in(in_reg_wire_7[203]),
    .out(out47)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1228]),
    .in(in_reg_wire_7[204]),
    .out(out51)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1229]),
    .in(in_reg_wire_7[205]),
    .out(out55)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1230]),
    .in(in_reg_wire_7[206]),
    .out(out59)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1231]),
    .in(in_reg_wire_7[207]),
    .out(out63)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1232]),
    .in(in_reg_wire_7[208]),
    .out(out67)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1233]),
    .in(in_reg_wire_7[209]),
    .out(out71)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1234]),
    .in(in_reg_wire_7[210]),
    .out(out75)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1235]),
    .in(in_reg_wire_7[211]),
    .out(out79)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1236]),
    .in(in_reg_wire_7[212]),
    .out(out83)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1237]),
    .in(in_reg_wire_7[213]),
    .out(out87)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1238]),
    .in(in_reg_wire_7[214]),
    .out(out91)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1239]),
    .in(in_reg_wire_7[215]),
    .out(out95)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1240]),
    .in(in_reg_wire_7[216]),
    .out(out99)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1241]),
    .in(in_reg_wire_7[217]),
    .out(out103)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1242]),
    .in(in_reg_wire_7[218]),
    .out(out107)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1243]),
    .in(in_reg_wire_7[219]),
    .out(out111)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1244]),
    .in(in_reg_wire_7[220]),
    .out(out115)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1245]),
    .in(in_reg_wire_7[221]),
    .out(out119)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1246]),
    .in(in_reg_wire_7[222]),
    .out(out123)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1247]),
    .in(in_reg_wire_7[223]),
    .out(out127)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1248]),
    .in(in_reg_wire_7[224]),
    .out(out131)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1249]),
    .in(in_reg_wire_7[225]),
    .out(out135)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1250]),
    .in(in_reg_wire_7[226]),
    .out(out139)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1251]),
    .in(in_reg_wire_7[227]),
    .out(out143)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1252]),
    .in(in_reg_wire_7[228]),
    .out(out147)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1253]),
    .in(in_reg_wire_7[229]),
    .out(out151)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1254]),
    .in(in_reg_wire_7[230]),
    .out(out155)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1255]),
    .in(in_reg_wire_7[231]),
    .out(out159)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1256]),
    .in(in_reg_wire_7[232]),
    .out(out163)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1257]),
    .in(in_reg_wire_7[233]),
    .out(out167)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1258]),
    .in(in_reg_wire_7[234]),
    .out(out171)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1259]),
    .in(in_reg_wire_7[235]),
    .out(out175)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1260]),
    .in(in_reg_wire_7[236]),
    .out(out179)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1261]),
    .in(in_reg_wire_7[237]),
    .out(out183)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1262]),
    .in(in_reg_wire_7[238]),
    .out(out187)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1263]),
    .in(in_reg_wire_7[239]),
    .out(out191)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1264]),
    .in(in_reg_wire_7[240]),
    .out(out195)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1265]),
    .in(in_reg_wire_7[241]),
    .out(out199)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1266]),
    .in(in_reg_wire_7[242]),
    .out(out203)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1267]),
    .in(in_reg_wire_7[243]),
    .out(out207)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1268]),
    .in(in_reg_wire_7[244]),
    .out(out211)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1269]),
    .in(in_reg_wire_7[245]),
    .out(out215)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1270]),
    .in(in_reg_wire_7[246]),
    .out(out219)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1271]),
    .in(in_reg_wire_7[247]),
    .out(out223)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1272]),
    .in(in_reg_wire_7[248]),
    .out(out227)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1273]),
    .in(in_reg_wire_7[249]),
    .out(out231)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1274]),
    .in(in_reg_wire_7[250]),
    .out(out235)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1275]),
    .in(in_reg_wire_7[251]),
    .out(out239)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1276]),
    .in(in_reg_wire_7[252]),
    .out(out243)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1277]),
    .in(in_reg_wire_7[253]),
    .out(out247)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1278]),
    .in(in_reg_wire_7[254]),
    .out(out251)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en[1279]),
    .in(in_reg_wire_7[255]),
    .out(out255)
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_0
  (
    .sel(conf_out[7:0]),
    .in0(in_reg_wire_0[0]),
    .in1(in_reg_wire_0[64]),
    .in2(in_reg_wire_0[128]),
    .in3(in_reg_wire_0[192]),
    .out0(in_reg_wire_1[0]),
    .out1(in_reg_wire_1[1]),
    .out2(in_reg_wire_1[2]),
    .out3(in_reg_wire_1[3])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_1
  (
    .sel(conf_out[15:8]),
    .in0(in_reg_wire_0[1]),
    .in1(in_reg_wire_0[65]),
    .in2(in_reg_wire_0[129]),
    .in3(in_reg_wire_0[193]),
    .out0(in_reg_wire_1[4]),
    .out1(in_reg_wire_1[5]),
    .out2(in_reg_wire_1[6]),
    .out3(in_reg_wire_1[7])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_2
  (
    .sel(conf_out[23:16]),
    .in0(in_reg_wire_0[2]),
    .in1(in_reg_wire_0[66]),
    .in2(in_reg_wire_0[130]),
    .in3(in_reg_wire_0[194]),
    .out0(in_reg_wire_1[8]),
    .out1(in_reg_wire_1[9]),
    .out2(in_reg_wire_1[10]),
    .out3(in_reg_wire_1[11])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_3
  (
    .sel(conf_out[31:24]),
    .in0(in_reg_wire_0[3]),
    .in1(in_reg_wire_0[67]),
    .in2(in_reg_wire_0[131]),
    .in3(in_reg_wire_0[195]),
    .out0(in_reg_wire_1[12]),
    .out1(in_reg_wire_1[13]),
    .out2(in_reg_wire_1[14]),
    .out3(in_reg_wire_1[15])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_4
  (
    .sel(conf_out[39:32]),
    .in0(in_reg_wire_0[4]),
    .in1(in_reg_wire_0[68]),
    .in2(in_reg_wire_0[132]),
    .in3(in_reg_wire_0[196]),
    .out0(in_reg_wire_1[16]),
    .out1(in_reg_wire_1[17]),
    .out2(in_reg_wire_1[18]),
    .out3(in_reg_wire_1[19])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_5
  (
    .sel(conf_out[47:40]),
    .in0(in_reg_wire_0[5]),
    .in1(in_reg_wire_0[69]),
    .in2(in_reg_wire_0[133]),
    .in3(in_reg_wire_0[197]),
    .out0(in_reg_wire_1[20]),
    .out1(in_reg_wire_1[21]),
    .out2(in_reg_wire_1[22]),
    .out3(in_reg_wire_1[23])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_6
  (
    .sel(conf_out[55:48]),
    .in0(in_reg_wire_0[6]),
    .in1(in_reg_wire_0[70]),
    .in2(in_reg_wire_0[134]),
    .in3(in_reg_wire_0[198]),
    .out0(in_reg_wire_1[24]),
    .out1(in_reg_wire_1[25]),
    .out2(in_reg_wire_1[26]),
    .out3(in_reg_wire_1[27])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_7
  (
    .sel(conf_out[63:56]),
    .in0(in_reg_wire_0[7]),
    .in1(in_reg_wire_0[71]),
    .in2(in_reg_wire_0[135]),
    .in3(in_reg_wire_0[199]),
    .out0(in_reg_wire_1[28]),
    .out1(in_reg_wire_1[29]),
    .out2(in_reg_wire_1[30]),
    .out3(in_reg_wire_1[31])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_8
  (
    .sel(conf_out[71:64]),
    .in0(in_reg_wire_0[8]),
    .in1(in_reg_wire_0[72]),
    .in2(in_reg_wire_0[136]),
    .in3(in_reg_wire_0[200]),
    .out0(in_reg_wire_1[32]),
    .out1(in_reg_wire_1[33]),
    .out2(in_reg_wire_1[34]),
    .out3(in_reg_wire_1[35])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_9
  (
    .sel(conf_out[79:72]),
    .in0(in_reg_wire_0[9]),
    .in1(in_reg_wire_0[73]),
    .in2(in_reg_wire_0[137]),
    .in3(in_reg_wire_0[201]),
    .out0(in_reg_wire_1[36]),
    .out1(in_reg_wire_1[37]),
    .out2(in_reg_wire_1[38]),
    .out3(in_reg_wire_1[39])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_10
  (
    .sel(conf_out[87:80]),
    .in0(in_reg_wire_0[10]),
    .in1(in_reg_wire_0[74]),
    .in2(in_reg_wire_0[138]),
    .in3(in_reg_wire_0[202]),
    .out0(in_reg_wire_1[40]),
    .out1(in_reg_wire_1[41]),
    .out2(in_reg_wire_1[42]),
    .out3(in_reg_wire_1[43])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_11
  (
    .sel(conf_out[95:88]),
    .in0(in_reg_wire_0[11]),
    .in1(in_reg_wire_0[75]),
    .in2(in_reg_wire_0[139]),
    .in3(in_reg_wire_0[203]),
    .out0(in_reg_wire_1[44]),
    .out1(in_reg_wire_1[45]),
    .out2(in_reg_wire_1[46]),
    .out3(in_reg_wire_1[47])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_12
  (
    .sel(conf_out[103:96]),
    .in0(in_reg_wire_0[12]),
    .in1(in_reg_wire_0[76]),
    .in2(in_reg_wire_0[140]),
    .in3(in_reg_wire_0[204]),
    .out0(in_reg_wire_1[48]),
    .out1(in_reg_wire_1[49]),
    .out2(in_reg_wire_1[50]),
    .out3(in_reg_wire_1[51])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_13
  (
    .sel(conf_out[111:104]),
    .in0(in_reg_wire_0[13]),
    .in1(in_reg_wire_0[77]),
    .in2(in_reg_wire_0[141]),
    .in3(in_reg_wire_0[205]),
    .out0(in_reg_wire_1[52]),
    .out1(in_reg_wire_1[53]),
    .out2(in_reg_wire_1[54]),
    .out3(in_reg_wire_1[55])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_14
  (
    .sel(conf_out[119:112]),
    .in0(in_reg_wire_0[14]),
    .in1(in_reg_wire_0[78]),
    .in2(in_reg_wire_0[142]),
    .in3(in_reg_wire_0[206]),
    .out0(in_reg_wire_1[56]),
    .out1(in_reg_wire_1[57]),
    .out2(in_reg_wire_1[58]),
    .out3(in_reg_wire_1[59])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_15
  (
    .sel(conf_out[127:120]),
    .in0(in_reg_wire_0[15]),
    .in1(in_reg_wire_0[79]),
    .in2(in_reg_wire_0[143]),
    .in3(in_reg_wire_0[207]),
    .out0(in_reg_wire_1[60]),
    .out1(in_reg_wire_1[61]),
    .out2(in_reg_wire_1[62]),
    .out3(in_reg_wire_1[63])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_16
  (
    .sel(conf_out[135:128]),
    .in0(in_reg_wire_0[16]),
    .in1(in_reg_wire_0[80]),
    .in2(in_reg_wire_0[144]),
    .in3(in_reg_wire_0[208]),
    .out0(in_reg_wire_1[64]),
    .out1(in_reg_wire_1[65]),
    .out2(in_reg_wire_1[66]),
    .out3(in_reg_wire_1[67])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_17
  (
    .sel(conf_out[143:136]),
    .in0(in_reg_wire_0[17]),
    .in1(in_reg_wire_0[81]),
    .in2(in_reg_wire_0[145]),
    .in3(in_reg_wire_0[209]),
    .out0(in_reg_wire_1[68]),
    .out1(in_reg_wire_1[69]),
    .out2(in_reg_wire_1[70]),
    .out3(in_reg_wire_1[71])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_18
  (
    .sel(conf_out[151:144]),
    .in0(in_reg_wire_0[18]),
    .in1(in_reg_wire_0[82]),
    .in2(in_reg_wire_0[146]),
    .in3(in_reg_wire_0[210]),
    .out0(in_reg_wire_1[72]),
    .out1(in_reg_wire_1[73]),
    .out2(in_reg_wire_1[74]),
    .out3(in_reg_wire_1[75])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_19
  (
    .sel(conf_out[159:152]),
    .in0(in_reg_wire_0[19]),
    .in1(in_reg_wire_0[83]),
    .in2(in_reg_wire_0[147]),
    .in3(in_reg_wire_0[211]),
    .out0(in_reg_wire_1[76]),
    .out1(in_reg_wire_1[77]),
    .out2(in_reg_wire_1[78]),
    .out3(in_reg_wire_1[79])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_20
  (
    .sel(conf_out[167:160]),
    .in0(in_reg_wire_0[20]),
    .in1(in_reg_wire_0[84]),
    .in2(in_reg_wire_0[148]),
    .in3(in_reg_wire_0[212]),
    .out0(in_reg_wire_1[80]),
    .out1(in_reg_wire_1[81]),
    .out2(in_reg_wire_1[82]),
    .out3(in_reg_wire_1[83])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_21
  (
    .sel(conf_out[175:168]),
    .in0(in_reg_wire_0[21]),
    .in1(in_reg_wire_0[85]),
    .in2(in_reg_wire_0[149]),
    .in3(in_reg_wire_0[213]),
    .out0(in_reg_wire_1[84]),
    .out1(in_reg_wire_1[85]),
    .out2(in_reg_wire_1[86]),
    .out3(in_reg_wire_1[87])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_22
  (
    .sel(conf_out[183:176]),
    .in0(in_reg_wire_0[22]),
    .in1(in_reg_wire_0[86]),
    .in2(in_reg_wire_0[150]),
    .in3(in_reg_wire_0[214]),
    .out0(in_reg_wire_1[88]),
    .out1(in_reg_wire_1[89]),
    .out2(in_reg_wire_1[90]),
    .out3(in_reg_wire_1[91])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_23
  (
    .sel(conf_out[191:184]),
    .in0(in_reg_wire_0[23]),
    .in1(in_reg_wire_0[87]),
    .in2(in_reg_wire_0[151]),
    .in3(in_reg_wire_0[215]),
    .out0(in_reg_wire_1[92]),
    .out1(in_reg_wire_1[93]),
    .out2(in_reg_wire_1[94]),
    .out3(in_reg_wire_1[95])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_24
  (
    .sel(conf_out[199:192]),
    .in0(in_reg_wire_0[24]),
    .in1(in_reg_wire_0[88]),
    .in2(in_reg_wire_0[152]),
    .in3(in_reg_wire_0[216]),
    .out0(in_reg_wire_1[96]),
    .out1(in_reg_wire_1[97]),
    .out2(in_reg_wire_1[98]),
    .out3(in_reg_wire_1[99])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_25
  (
    .sel(conf_out[207:200]),
    .in0(in_reg_wire_0[25]),
    .in1(in_reg_wire_0[89]),
    .in2(in_reg_wire_0[153]),
    .in3(in_reg_wire_0[217]),
    .out0(in_reg_wire_1[100]),
    .out1(in_reg_wire_1[101]),
    .out2(in_reg_wire_1[102]),
    .out3(in_reg_wire_1[103])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_26
  (
    .sel(conf_out[215:208]),
    .in0(in_reg_wire_0[26]),
    .in1(in_reg_wire_0[90]),
    .in2(in_reg_wire_0[154]),
    .in3(in_reg_wire_0[218]),
    .out0(in_reg_wire_1[104]),
    .out1(in_reg_wire_1[105]),
    .out2(in_reg_wire_1[106]),
    .out3(in_reg_wire_1[107])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_27
  (
    .sel(conf_out[223:216]),
    .in0(in_reg_wire_0[27]),
    .in1(in_reg_wire_0[91]),
    .in2(in_reg_wire_0[155]),
    .in3(in_reg_wire_0[219]),
    .out0(in_reg_wire_1[108]),
    .out1(in_reg_wire_1[109]),
    .out2(in_reg_wire_1[110]),
    .out3(in_reg_wire_1[111])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_28
  (
    .sel(conf_out[231:224]),
    .in0(in_reg_wire_0[28]),
    .in1(in_reg_wire_0[92]),
    .in2(in_reg_wire_0[156]),
    .in3(in_reg_wire_0[220]),
    .out0(in_reg_wire_1[112]),
    .out1(in_reg_wire_1[113]),
    .out2(in_reg_wire_1[114]),
    .out3(in_reg_wire_1[115])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_29
  (
    .sel(conf_out[239:232]),
    .in0(in_reg_wire_0[29]),
    .in1(in_reg_wire_0[93]),
    .in2(in_reg_wire_0[157]),
    .in3(in_reg_wire_0[221]),
    .out0(in_reg_wire_1[116]),
    .out1(in_reg_wire_1[117]),
    .out2(in_reg_wire_1[118]),
    .out3(in_reg_wire_1[119])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_30
  (
    .sel(conf_out[247:240]),
    .in0(in_reg_wire_0[30]),
    .in1(in_reg_wire_0[94]),
    .in2(in_reg_wire_0[158]),
    .in3(in_reg_wire_0[222]),
    .out0(in_reg_wire_1[120]),
    .out1(in_reg_wire_1[121]),
    .out2(in_reg_wire_1[122]),
    .out3(in_reg_wire_1[123])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_31
  (
    .sel(conf_out[255:248]),
    .in0(in_reg_wire_0[31]),
    .in1(in_reg_wire_0[95]),
    .in2(in_reg_wire_0[159]),
    .in3(in_reg_wire_0[223]),
    .out0(in_reg_wire_1[124]),
    .out1(in_reg_wire_1[125]),
    .out2(in_reg_wire_1[126]),
    .out3(in_reg_wire_1[127])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_32
  (
    .sel(conf_out[263:256]),
    .in0(in_reg_wire_0[32]),
    .in1(in_reg_wire_0[96]),
    .in2(in_reg_wire_0[160]),
    .in3(in_reg_wire_0[224]),
    .out0(in_reg_wire_1[128]),
    .out1(in_reg_wire_1[129]),
    .out2(in_reg_wire_1[130]),
    .out3(in_reg_wire_1[131])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_33
  (
    .sel(conf_out[271:264]),
    .in0(in_reg_wire_0[33]),
    .in1(in_reg_wire_0[97]),
    .in2(in_reg_wire_0[161]),
    .in3(in_reg_wire_0[225]),
    .out0(in_reg_wire_1[132]),
    .out1(in_reg_wire_1[133]),
    .out2(in_reg_wire_1[134]),
    .out3(in_reg_wire_1[135])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_34
  (
    .sel(conf_out[279:272]),
    .in0(in_reg_wire_0[34]),
    .in1(in_reg_wire_0[98]),
    .in2(in_reg_wire_0[162]),
    .in3(in_reg_wire_0[226]),
    .out0(in_reg_wire_1[136]),
    .out1(in_reg_wire_1[137]),
    .out2(in_reg_wire_1[138]),
    .out3(in_reg_wire_1[139])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_35
  (
    .sel(conf_out[287:280]),
    .in0(in_reg_wire_0[35]),
    .in1(in_reg_wire_0[99]),
    .in2(in_reg_wire_0[163]),
    .in3(in_reg_wire_0[227]),
    .out0(in_reg_wire_1[140]),
    .out1(in_reg_wire_1[141]),
    .out2(in_reg_wire_1[142]),
    .out3(in_reg_wire_1[143])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_36
  (
    .sel(conf_out[295:288]),
    .in0(in_reg_wire_0[36]),
    .in1(in_reg_wire_0[100]),
    .in2(in_reg_wire_0[164]),
    .in3(in_reg_wire_0[228]),
    .out0(in_reg_wire_1[144]),
    .out1(in_reg_wire_1[145]),
    .out2(in_reg_wire_1[146]),
    .out3(in_reg_wire_1[147])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_37
  (
    .sel(conf_out[303:296]),
    .in0(in_reg_wire_0[37]),
    .in1(in_reg_wire_0[101]),
    .in2(in_reg_wire_0[165]),
    .in3(in_reg_wire_0[229]),
    .out0(in_reg_wire_1[148]),
    .out1(in_reg_wire_1[149]),
    .out2(in_reg_wire_1[150]),
    .out3(in_reg_wire_1[151])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_38
  (
    .sel(conf_out[311:304]),
    .in0(in_reg_wire_0[38]),
    .in1(in_reg_wire_0[102]),
    .in2(in_reg_wire_0[166]),
    .in3(in_reg_wire_0[230]),
    .out0(in_reg_wire_1[152]),
    .out1(in_reg_wire_1[153]),
    .out2(in_reg_wire_1[154]),
    .out3(in_reg_wire_1[155])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_39
  (
    .sel(conf_out[319:312]),
    .in0(in_reg_wire_0[39]),
    .in1(in_reg_wire_0[103]),
    .in2(in_reg_wire_0[167]),
    .in3(in_reg_wire_0[231]),
    .out0(in_reg_wire_1[156]),
    .out1(in_reg_wire_1[157]),
    .out2(in_reg_wire_1[158]),
    .out3(in_reg_wire_1[159])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_40
  (
    .sel(conf_out[327:320]),
    .in0(in_reg_wire_0[40]),
    .in1(in_reg_wire_0[104]),
    .in2(in_reg_wire_0[168]),
    .in3(in_reg_wire_0[232]),
    .out0(in_reg_wire_1[160]),
    .out1(in_reg_wire_1[161]),
    .out2(in_reg_wire_1[162]),
    .out3(in_reg_wire_1[163])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_41
  (
    .sel(conf_out[335:328]),
    .in0(in_reg_wire_0[41]),
    .in1(in_reg_wire_0[105]),
    .in2(in_reg_wire_0[169]),
    .in3(in_reg_wire_0[233]),
    .out0(in_reg_wire_1[164]),
    .out1(in_reg_wire_1[165]),
    .out2(in_reg_wire_1[166]),
    .out3(in_reg_wire_1[167])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_42
  (
    .sel(conf_out[343:336]),
    .in0(in_reg_wire_0[42]),
    .in1(in_reg_wire_0[106]),
    .in2(in_reg_wire_0[170]),
    .in3(in_reg_wire_0[234]),
    .out0(in_reg_wire_1[168]),
    .out1(in_reg_wire_1[169]),
    .out2(in_reg_wire_1[170]),
    .out3(in_reg_wire_1[171])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_43
  (
    .sel(conf_out[351:344]),
    .in0(in_reg_wire_0[43]),
    .in1(in_reg_wire_0[107]),
    .in2(in_reg_wire_0[171]),
    .in3(in_reg_wire_0[235]),
    .out0(in_reg_wire_1[172]),
    .out1(in_reg_wire_1[173]),
    .out2(in_reg_wire_1[174]),
    .out3(in_reg_wire_1[175])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_44
  (
    .sel(conf_out[359:352]),
    .in0(in_reg_wire_0[44]),
    .in1(in_reg_wire_0[108]),
    .in2(in_reg_wire_0[172]),
    .in3(in_reg_wire_0[236]),
    .out0(in_reg_wire_1[176]),
    .out1(in_reg_wire_1[177]),
    .out2(in_reg_wire_1[178]),
    .out3(in_reg_wire_1[179])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_45
  (
    .sel(conf_out[367:360]),
    .in0(in_reg_wire_0[45]),
    .in1(in_reg_wire_0[109]),
    .in2(in_reg_wire_0[173]),
    .in3(in_reg_wire_0[237]),
    .out0(in_reg_wire_1[180]),
    .out1(in_reg_wire_1[181]),
    .out2(in_reg_wire_1[182]),
    .out3(in_reg_wire_1[183])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_46
  (
    .sel(conf_out[375:368]),
    .in0(in_reg_wire_0[46]),
    .in1(in_reg_wire_0[110]),
    .in2(in_reg_wire_0[174]),
    .in3(in_reg_wire_0[238]),
    .out0(in_reg_wire_1[184]),
    .out1(in_reg_wire_1[185]),
    .out2(in_reg_wire_1[186]),
    .out3(in_reg_wire_1[187])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_47
  (
    .sel(conf_out[383:376]),
    .in0(in_reg_wire_0[47]),
    .in1(in_reg_wire_0[111]),
    .in2(in_reg_wire_0[175]),
    .in3(in_reg_wire_0[239]),
    .out0(in_reg_wire_1[188]),
    .out1(in_reg_wire_1[189]),
    .out2(in_reg_wire_1[190]),
    .out3(in_reg_wire_1[191])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_48
  (
    .sel(conf_out[391:384]),
    .in0(in_reg_wire_0[48]),
    .in1(in_reg_wire_0[112]),
    .in2(in_reg_wire_0[176]),
    .in3(in_reg_wire_0[240]),
    .out0(in_reg_wire_1[192]),
    .out1(in_reg_wire_1[193]),
    .out2(in_reg_wire_1[194]),
    .out3(in_reg_wire_1[195])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_49
  (
    .sel(conf_out[399:392]),
    .in0(in_reg_wire_0[49]),
    .in1(in_reg_wire_0[113]),
    .in2(in_reg_wire_0[177]),
    .in3(in_reg_wire_0[241]),
    .out0(in_reg_wire_1[196]),
    .out1(in_reg_wire_1[197]),
    .out2(in_reg_wire_1[198]),
    .out3(in_reg_wire_1[199])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_50
  (
    .sel(conf_out[407:400]),
    .in0(in_reg_wire_0[50]),
    .in1(in_reg_wire_0[114]),
    .in2(in_reg_wire_0[178]),
    .in3(in_reg_wire_0[242]),
    .out0(in_reg_wire_1[200]),
    .out1(in_reg_wire_1[201]),
    .out2(in_reg_wire_1[202]),
    .out3(in_reg_wire_1[203])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_51
  (
    .sel(conf_out[415:408]),
    .in0(in_reg_wire_0[51]),
    .in1(in_reg_wire_0[115]),
    .in2(in_reg_wire_0[179]),
    .in3(in_reg_wire_0[243]),
    .out0(in_reg_wire_1[204]),
    .out1(in_reg_wire_1[205]),
    .out2(in_reg_wire_1[206]),
    .out3(in_reg_wire_1[207])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_52
  (
    .sel(conf_out[423:416]),
    .in0(in_reg_wire_0[52]),
    .in1(in_reg_wire_0[116]),
    .in2(in_reg_wire_0[180]),
    .in3(in_reg_wire_0[244]),
    .out0(in_reg_wire_1[208]),
    .out1(in_reg_wire_1[209]),
    .out2(in_reg_wire_1[210]),
    .out3(in_reg_wire_1[211])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_53
  (
    .sel(conf_out[431:424]),
    .in0(in_reg_wire_0[53]),
    .in1(in_reg_wire_0[117]),
    .in2(in_reg_wire_0[181]),
    .in3(in_reg_wire_0[245]),
    .out0(in_reg_wire_1[212]),
    .out1(in_reg_wire_1[213]),
    .out2(in_reg_wire_1[214]),
    .out3(in_reg_wire_1[215])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_54
  (
    .sel(conf_out[439:432]),
    .in0(in_reg_wire_0[54]),
    .in1(in_reg_wire_0[118]),
    .in2(in_reg_wire_0[182]),
    .in3(in_reg_wire_0[246]),
    .out0(in_reg_wire_1[216]),
    .out1(in_reg_wire_1[217]),
    .out2(in_reg_wire_1[218]),
    .out3(in_reg_wire_1[219])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_55
  (
    .sel(conf_out[447:440]),
    .in0(in_reg_wire_0[55]),
    .in1(in_reg_wire_0[119]),
    .in2(in_reg_wire_0[183]),
    .in3(in_reg_wire_0[247]),
    .out0(in_reg_wire_1[220]),
    .out1(in_reg_wire_1[221]),
    .out2(in_reg_wire_1[222]),
    .out3(in_reg_wire_1[223])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_56
  (
    .sel(conf_out[455:448]),
    .in0(in_reg_wire_0[56]),
    .in1(in_reg_wire_0[120]),
    .in2(in_reg_wire_0[184]),
    .in3(in_reg_wire_0[248]),
    .out0(in_reg_wire_1[224]),
    .out1(in_reg_wire_1[225]),
    .out2(in_reg_wire_1[226]),
    .out3(in_reg_wire_1[227])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_57
  (
    .sel(conf_out[463:456]),
    .in0(in_reg_wire_0[57]),
    .in1(in_reg_wire_0[121]),
    .in2(in_reg_wire_0[185]),
    .in3(in_reg_wire_0[249]),
    .out0(in_reg_wire_1[228]),
    .out1(in_reg_wire_1[229]),
    .out2(in_reg_wire_1[230]),
    .out3(in_reg_wire_1[231])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_58
  (
    .sel(conf_out[471:464]),
    .in0(in_reg_wire_0[58]),
    .in1(in_reg_wire_0[122]),
    .in2(in_reg_wire_0[186]),
    .in3(in_reg_wire_0[250]),
    .out0(in_reg_wire_1[232]),
    .out1(in_reg_wire_1[233]),
    .out2(in_reg_wire_1[234]),
    .out3(in_reg_wire_1[235])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_59
  (
    .sel(conf_out[479:472]),
    .in0(in_reg_wire_0[59]),
    .in1(in_reg_wire_0[123]),
    .in2(in_reg_wire_0[187]),
    .in3(in_reg_wire_0[251]),
    .out0(in_reg_wire_1[236]),
    .out1(in_reg_wire_1[237]),
    .out2(in_reg_wire_1[238]),
    .out3(in_reg_wire_1[239])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_60
  (
    .sel(conf_out[487:480]),
    .in0(in_reg_wire_0[60]),
    .in1(in_reg_wire_0[124]),
    .in2(in_reg_wire_0[188]),
    .in3(in_reg_wire_0[252]),
    .out0(in_reg_wire_1[240]),
    .out1(in_reg_wire_1[241]),
    .out2(in_reg_wire_1[242]),
    .out3(in_reg_wire_1[243])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_61
  (
    .sel(conf_out[495:488]),
    .in0(in_reg_wire_0[61]),
    .in1(in_reg_wire_0[125]),
    .in2(in_reg_wire_0[189]),
    .in3(in_reg_wire_0[253]),
    .out0(in_reg_wire_1[244]),
    .out1(in_reg_wire_1[245]),
    .out2(in_reg_wire_1[246]),
    .out3(in_reg_wire_1[247])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_62
  (
    .sel(conf_out[503:496]),
    .in0(in_reg_wire_0[62]),
    .in1(in_reg_wire_0[126]),
    .in2(in_reg_wire_0[190]),
    .in3(in_reg_wire_0[254]),
    .out0(in_reg_wire_1[248]),
    .out1(in_reg_wire_1[249]),
    .out2(in_reg_wire_1[250]),
    .out3(in_reg_wire_1[251])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_0_63
  (
    .sel(conf_out[511:504]),
    .in0(in_reg_wire_0[63]),
    .in1(in_reg_wire_0[127]),
    .in2(in_reg_wire_0[191]),
    .in3(in_reg_wire_0[255]),
    .out0(in_reg_wire_1[252]),
    .out1(in_reg_wire_1[253]),
    .out2(in_reg_wire_1[254]),
    .out3(in_reg_wire_1[255])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_0
  (
    .sel(conf_out[519:512]),
    .in0(in_reg_wire_2[0]),
    .in1(in_reg_wire_2[64]),
    .in2(in_reg_wire_2[128]),
    .in3(in_reg_wire_2[192]),
    .out0(in_reg_wire_3[0]),
    .out1(in_reg_wire_3[1]),
    .out2(in_reg_wire_3[2]),
    .out3(in_reg_wire_3[3])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_1
  (
    .sel(conf_out[527:520]),
    .in0(in_reg_wire_2[1]),
    .in1(in_reg_wire_2[65]),
    .in2(in_reg_wire_2[129]),
    .in3(in_reg_wire_2[193]),
    .out0(in_reg_wire_3[4]),
    .out1(in_reg_wire_3[5]),
    .out2(in_reg_wire_3[6]),
    .out3(in_reg_wire_3[7])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_2
  (
    .sel(conf_out[535:528]),
    .in0(in_reg_wire_2[2]),
    .in1(in_reg_wire_2[66]),
    .in2(in_reg_wire_2[130]),
    .in3(in_reg_wire_2[194]),
    .out0(in_reg_wire_3[8]),
    .out1(in_reg_wire_3[9]),
    .out2(in_reg_wire_3[10]),
    .out3(in_reg_wire_3[11])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_3
  (
    .sel(conf_out[543:536]),
    .in0(in_reg_wire_2[3]),
    .in1(in_reg_wire_2[67]),
    .in2(in_reg_wire_2[131]),
    .in3(in_reg_wire_2[195]),
    .out0(in_reg_wire_3[12]),
    .out1(in_reg_wire_3[13]),
    .out2(in_reg_wire_3[14]),
    .out3(in_reg_wire_3[15])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_4
  (
    .sel(conf_out[551:544]),
    .in0(in_reg_wire_2[4]),
    .in1(in_reg_wire_2[68]),
    .in2(in_reg_wire_2[132]),
    .in3(in_reg_wire_2[196]),
    .out0(in_reg_wire_3[16]),
    .out1(in_reg_wire_3[17]),
    .out2(in_reg_wire_3[18]),
    .out3(in_reg_wire_3[19])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_5
  (
    .sel(conf_out[559:552]),
    .in0(in_reg_wire_2[5]),
    .in1(in_reg_wire_2[69]),
    .in2(in_reg_wire_2[133]),
    .in3(in_reg_wire_2[197]),
    .out0(in_reg_wire_3[20]),
    .out1(in_reg_wire_3[21]),
    .out2(in_reg_wire_3[22]),
    .out3(in_reg_wire_3[23])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_6
  (
    .sel(conf_out[567:560]),
    .in0(in_reg_wire_2[6]),
    .in1(in_reg_wire_2[70]),
    .in2(in_reg_wire_2[134]),
    .in3(in_reg_wire_2[198]),
    .out0(in_reg_wire_3[24]),
    .out1(in_reg_wire_3[25]),
    .out2(in_reg_wire_3[26]),
    .out3(in_reg_wire_3[27])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_7
  (
    .sel(conf_out[575:568]),
    .in0(in_reg_wire_2[7]),
    .in1(in_reg_wire_2[71]),
    .in2(in_reg_wire_2[135]),
    .in3(in_reg_wire_2[199]),
    .out0(in_reg_wire_3[28]),
    .out1(in_reg_wire_3[29]),
    .out2(in_reg_wire_3[30]),
    .out3(in_reg_wire_3[31])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_8
  (
    .sel(conf_out[583:576]),
    .in0(in_reg_wire_2[8]),
    .in1(in_reg_wire_2[72]),
    .in2(in_reg_wire_2[136]),
    .in3(in_reg_wire_2[200]),
    .out0(in_reg_wire_3[32]),
    .out1(in_reg_wire_3[33]),
    .out2(in_reg_wire_3[34]),
    .out3(in_reg_wire_3[35])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_9
  (
    .sel(conf_out[591:584]),
    .in0(in_reg_wire_2[9]),
    .in1(in_reg_wire_2[73]),
    .in2(in_reg_wire_2[137]),
    .in3(in_reg_wire_2[201]),
    .out0(in_reg_wire_3[36]),
    .out1(in_reg_wire_3[37]),
    .out2(in_reg_wire_3[38]),
    .out3(in_reg_wire_3[39])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_10
  (
    .sel(conf_out[599:592]),
    .in0(in_reg_wire_2[10]),
    .in1(in_reg_wire_2[74]),
    .in2(in_reg_wire_2[138]),
    .in3(in_reg_wire_2[202]),
    .out0(in_reg_wire_3[40]),
    .out1(in_reg_wire_3[41]),
    .out2(in_reg_wire_3[42]),
    .out3(in_reg_wire_3[43])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_11
  (
    .sel(conf_out[607:600]),
    .in0(in_reg_wire_2[11]),
    .in1(in_reg_wire_2[75]),
    .in2(in_reg_wire_2[139]),
    .in3(in_reg_wire_2[203]),
    .out0(in_reg_wire_3[44]),
    .out1(in_reg_wire_3[45]),
    .out2(in_reg_wire_3[46]),
    .out3(in_reg_wire_3[47])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_12
  (
    .sel(conf_out[615:608]),
    .in0(in_reg_wire_2[12]),
    .in1(in_reg_wire_2[76]),
    .in2(in_reg_wire_2[140]),
    .in3(in_reg_wire_2[204]),
    .out0(in_reg_wire_3[48]),
    .out1(in_reg_wire_3[49]),
    .out2(in_reg_wire_3[50]),
    .out3(in_reg_wire_3[51])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_13
  (
    .sel(conf_out[623:616]),
    .in0(in_reg_wire_2[13]),
    .in1(in_reg_wire_2[77]),
    .in2(in_reg_wire_2[141]),
    .in3(in_reg_wire_2[205]),
    .out0(in_reg_wire_3[52]),
    .out1(in_reg_wire_3[53]),
    .out2(in_reg_wire_3[54]),
    .out3(in_reg_wire_3[55])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_14
  (
    .sel(conf_out[631:624]),
    .in0(in_reg_wire_2[14]),
    .in1(in_reg_wire_2[78]),
    .in2(in_reg_wire_2[142]),
    .in3(in_reg_wire_2[206]),
    .out0(in_reg_wire_3[56]),
    .out1(in_reg_wire_3[57]),
    .out2(in_reg_wire_3[58]),
    .out3(in_reg_wire_3[59])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_15
  (
    .sel(conf_out[639:632]),
    .in0(in_reg_wire_2[15]),
    .in1(in_reg_wire_2[79]),
    .in2(in_reg_wire_2[143]),
    .in3(in_reg_wire_2[207]),
    .out0(in_reg_wire_3[60]),
    .out1(in_reg_wire_3[61]),
    .out2(in_reg_wire_3[62]),
    .out3(in_reg_wire_3[63])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_16
  (
    .sel(conf_out[647:640]),
    .in0(in_reg_wire_2[16]),
    .in1(in_reg_wire_2[80]),
    .in2(in_reg_wire_2[144]),
    .in3(in_reg_wire_2[208]),
    .out0(in_reg_wire_3[64]),
    .out1(in_reg_wire_3[65]),
    .out2(in_reg_wire_3[66]),
    .out3(in_reg_wire_3[67])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_17
  (
    .sel(conf_out[655:648]),
    .in0(in_reg_wire_2[17]),
    .in1(in_reg_wire_2[81]),
    .in2(in_reg_wire_2[145]),
    .in3(in_reg_wire_2[209]),
    .out0(in_reg_wire_3[68]),
    .out1(in_reg_wire_3[69]),
    .out2(in_reg_wire_3[70]),
    .out3(in_reg_wire_3[71])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_18
  (
    .sel(conf_out[663:656]),
    .in0(in_reg_wire_2[18]),
    .in1(in_reg_wire_2[82]),
    .in2(in_reg_wire_2[146]),
    .in3(in_reg_wire_2[210]),
    .out0(in_reg_wire_3[72]),
    .out1(in_reg_wire_3[73]),
    .out2(in_reg_wire_3[74]),
    .out3(in_reg_wire_3[75])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_19
  (
    .sel(conf_out[671:664]),
    .in0(in_reg_wire_2[19]),
    .in1(in_reg_wire_2[83]),
    .in2(in_reg_wire_2[147]),
    .in3(in_reg_wire_2[211]),
    .out0(in_reg_wire_3[76]),
    .out1(in_reg_wire_3[77]),
    .out2(in_reg_wire_3[78]),
    .out3(in_reg_wire_3[79])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_20
  (
    .sel(conf_out[679:672]),
    .in0(in_reg_wire_2[20]),
    .in1(in_reg_wire_2[84]),
    .in2(in_reg_wire_2[148]),
    .in3(in_reg_wire_2[212]),
    .out0(in_reg_wire_3[80]),
    .out1(in_reg_wire_3[81]),
    .out2(in_reg_wire_3[82]),
    .out3(in_reg_wire_3[83])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_21
  (
    .sel(conf_out[687:680]),
    .in0(in_reg_wire_2[21]),
    .in1(in_reg_wire_2[85]),
    .in2(in_reg_wire_2[149]),
    .in3(in_reg_wire_2[213]),
    .out0(in_reg_wire_3[84]),
    .out1(in_reg_wire_3[85]),
    .out2(in_reg_wire_3[86]),
    .out3(in_reg_wire_3[87])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_22
  (
    .sel(conf_out[695:688]),
    .in0(in_reg_wire_2[22]),
    .in1(in_reg_wire_2[86]),
    .in2(in_reg_wire_2[150]),
    .in3(in_reg_wire_2[214]),
    .out0(in_reg_wire_3[88]),
    .out1(in_reg_wire_3[89]),
    .out2(in_reg_wire_3[90]),
    .out3(in_reg_wire_3[91])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_23
  (
    .sel(conf_out[703:696]),
    .in0(in_reg_wire_2[23]),
    .in1(in_reg_wire_2[87]),
    .in2(in_reg_wire_2[151]),
    .in3(in_reg_wire_2[215]),
    .out0(in_reg_wire_3[92]),
    .out1(in_reg_wire_3[93]),
    .out2(in_reg_wire_3[94]),
    .out3(in_reg_wire_3[95])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_24
  (
    .sel(conf_out[711:704]),
    .in0(in_reg_wire_2[24]),
    .in1(in_reg_wire_2[88]),
    .in2(in_reg_wire_2[152]),
    .in3(in_reg_wire_2[216]),
    .out0(in_reg_wire_3[96]),
    .out1(in_reg_wire_3[97]),
    .out2(in_reg_wire_3[98]),
    .out3(in_reg_wire_3[99])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_25
  (
    .sel(conf_out[719:712]),
    .in0(in_reg_wire_2[25]),
    .in1(in_reg_wire_2[89]),
    .in2(in_reg_wire_2[153]),
    .in3(in_reg_wire_2[217]),
    .out0(in_reg_wire_3[100]),
    .out1(in_reg_wire_3[101]),
    .out2(in_reg_wire_3[102]),
    .out3(in_reg_wire_3[103])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_26
  (
    .sel(conf_out[727:720]),
    .in0(in_reg_wire_2[26]),
    .in1(in_reg_wire_2[90]),
    .in2(in_reg_wire_2[154]),
    .in3(in_reg_wire_2[218]),
    .out0(in_reg_wire_3[104]),
    .out1(in_reg_wire_3[105]),
    .out2(in_reg_wire_3[106]),
    .out3(in_reg_wire_3[107])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_27
  (
    .sel(conf_out[735:728]),
    .in0(in_reg_wire_2[27]),
    .in1(in_reg_wire_2[91]),
    .in2(in_reg_wire_2[155]),
    .in3(in_reg_wire_2[219]),
    .out0(in_reg_wire_3[108]),
    .out1(in_reg_wire_3[109]),
    .out2(in_reg_wire_3[110]),
    .out3(in_reg_wire_3[111])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_28
  (
    .sel(conf_out[743:736]),
    .in0(in_reg_wire_2[28]),
    .in1(in_reg_wire_2[92]),
    .in2(in_reg_wire_2[156]),
    .in3(in_reg_wire_2[220]),
    .out0(in_reg_wire_3[112]),
    .out1(in_reg_wire_3[113]),
    .out2(in_reg_wire_3[114]),
    .out3(in_reg_wire_3[115])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_29
  (
    .sel(conf_out[751:744]),
    .in0(in_reg_wire_2[29]),
    .in1(in_reg_wire_2[93]),
    .in2(in_reg_wire_2[157]),
    .in3(in_reg_wire_2[221]),
    .out0(in_reg_wire_3[116]),
    .out1(in_reg_wire_3[117]),
    .out2(in_reg_wire_3[118]),
    .out3(in_reg_wire_3[119])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_30
  (
    .sel(conf_out[759:752]),
    .in0(in_reg_wire_2[30]),
    .in1(in_reg_wire_2[94]),
    .in2(in_reg_wire_2[158]),
    .in3(in_reg_wire_2[222]),
    .out0(in_reg_wire_3[120]),
    .out1(in_reg_wire_3[121]),
    .out2(in_reg_wire_3[122]),
    .out3(in_reg_wire_3[123])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_31
  (
    .sel(conf_out[767:760]),
    .in0(in_reg_wire_2[31]),
    .in1(in_reg_wire_2[95]),
    .in2(in_reg_wire_2[159]),
    .in3(in_reg_wire_2[223]),
    .out0(in_reg_wire_3[124]),
    .out1(in_reg_wire_3[125]),
    .out2(in_reg_wire_3[126]),
    .out3(in_reg_wire_3[127])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_32
  (
    .sel(conf_out[775:768]),
    .in0(in_reg_wire_2[32]),
    .in1(in_reg_wire_2[96]),
    .in2(in_reg_wire_2[160]),
    .in3(in_reg_wire_2[224]),
    .out0(in_reg_wire_3[128]),
    .out1(in_reg_wire_3[129]),
    .out2(in_reg_wire_3[130]),
    .out3(in_reg_wire_3[131])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_33
  (
    .sel(conf_out[783:776]),
    .in0(in_reg_wire_2[33]),
    .in1(in_reg_wire_2[97]),
    .in2(in_reg_wire_2[161]),
    .in3(in_reg_wire_2[225]),
    .out0(in_reg_wire_3[132]),
    .out1(in_reg_wire_3[133]),
    .out2(in_reg_wire_3[134]),
    .out3(in_reg_wire_3[135])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_34
  (
    .sel(conf_out[791:784]),
    .in0(in_reg_wire_2[34]),
    .in1(in_reg_wire_2[98]),
    .in2(in_reg_wire_2[162]),
    .in3(in_reg_wire_2[226]),
    .out0(in_reg_wire_3[136]),
    .out1(in_reg_wire_3[137]),
    .out2(in_reg_wire_3[138]),
    .out3(in_reg_wire_3[139])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_35
  (
    .sel(conf_out[799:792]),
    .in0(in_reg_wire_2[35]),
    .in1(in_reg_wire_2[99]),
    .in2(in_reg_wire_2[163]),
    .in3(in_reg_wire_2[227]),
    .out0(in_reg_wire_3[140]),
    .out1(in_reg_wire_3[141]),
    .out2(in_reg_wire_3[142]),
    .out3(in_reg_wire_3[143])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_36
  (
    .sel(conf_out[807:800]),
    .in0(in_reg_wire_2[36]),
    .in1(in_reg_wire_2[100]),
    .in2(in_reg_wire_2[164]),
    .in3(in_reg_wire_2[228]),
    .out0(in_reg_wire_3[144]),
    .out1(in_reg_wire_3[145]),
    .out2(in_reg_wire_3[146]),
    .out3(in_reg_wire_3[147])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_37
  (
    .sel(conf_out[815:808]),
    .in0(in_reg_wire_2[37]),
    .in1(in_reg_wire_2[101]),
    .in2(in_reg_wire_2[165]),
    .in3(in_reg_wire_2[229]),
    .out0(in_reg_wire_3[148]),
    .out1(in_reg_wire_3[149]),
    .out2(in_reg_wire_3[150]),
    .out3(in_reg_wire_3[151])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_38
  (
    .sel(conf_out[823:816]),
    .in0(in_reg_wire_2[38]),
    .in1(in_reg_wire_2[102]),
    .in2(in_reg_wire_2[166]),
    .in3(in_reg_wire_2[230]),
    .out0(in_reg_wire_3[152]),
    .out1(in_reg_wire_3[153]),
    .out2(in_reg_wire_3[154]),
    .out3(in_reg_wire_3[155])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_39
  (
    .sel(conf_out[831:824]),
    .in0(in_reg_wire_2[39]),
    .in1(in_reg_wire_2[103]),
    .in2(in_reg_wire_2[167]),
    .in3(in_reg_wire_2[231]),
    .out0(in_reg_wire_3[156]),
    .out1(in_reg_wire_3[157]),
    .out2(in_reg_wire_3[158]),
    .out3(in_reg_wire_3[159])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_40
  (
    .sel(conf_out[839:832]),
    .in0(in_reg_wire_2[40]),
    .in1(in_reg_wire_2[104]),
    .in2(in_reg_wire_2[168]),
    .in3(in_reg_wire_2[232]),
    .out0(in_reg_wire_3[160]),
    .out1(in_reg_wire_3[161]),
    .out2(in_reg_wire_3[162]),
    .out3(in_reg_wire_3[163])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_41
  (
    .sel(conf_out[847:840]),
    .in0(in_reg_wire_2[41]),
    .in1(in_reg_wire_2[105]),
    .in2(in_reg_wire_2[169]),
    .in3(in_reg_wire_2[233]),
    .out0(in_reg_wire_3[164]),
    .out1(in_reg_wire_3[165]),
    .out2(in_reg_wire_3[166]),
    .out3(in_reg_wire_3[167])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_42
  (
    .sel(conf_out[855:848]),
    .in0(in_reg_wire_2[42]),
    .in1(in_reg_wire_2[106]),
    .in2(in_reg_wire_2[170]),
    .in3(in_reg_wire_2[234]),
    .out0(in_reg_wire_3[168]),
    .out1(in_reg_wire_3[169]),
    .out2(in_reg_wire_3[170]),
    .out3(in_reg_wire_3[171])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_43
  (
    .sel(conf_out[863:856]),
    .in0(in_reg_wire_2[43]),
    .in1(in_reg_wire_2[107]),
    .in2(in_reg_wire_2[171]),
    .in3(in_reg_wire_2[235]),
    .out0(in_reg_wire_3[172]),
    .out1(in_reg_wire_3[173]),
    .out2(in_reg_wire_3[174]),
    .out3(in_reg_wire_3[175])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_44
  (
    .sel(conf_out[871:864]),
    .in0(in_reg_wire_2[44]),
    .in1(in_reg_wire_2[108]),
    .in2(in_reg_wire_2[172]),
    .in3(in_reg_wire_2[236]),
    .out0(in_reg_wire_3[176]),
    .out1(in_reg_wire_3[177]),
    .out2(in_reg_wire_3[178]),
    .out3(in_reg_wire_3[179])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_45
  (
    .sel(conf_out[879:872]),
    .in0(in_reg_wire_2[45]),
    .in1(in_reg_wire_2[109]),
    .in2(in_reg_wire_2[173]),
    .in3(in_reg_wire_2[237]),
    .out0(in_reg_wire_3[180]),
    .out1(in_reg_wire_3[181]),
    .out2(in_reg_wire_3[182]),
    .out3(in_reg_wire_3[183])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_46
  (
    .sel(conf_out[887:880]),
    .in0(in_reg_wire_2[46]),
    .in1(in_reg_wire_2[110]),
    .in2(in_reg_wire_2[174]),
    .in3(in_reg_wire_2[238]),
    .out0(in_reg_wire_3[184]),
    .out1(in_reg_wire_3[185]),
    .out2(in_reg_wire_3[186]),
    .out3(in_reg_wire_3[187])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_47
  (
    .sel(conf_out[895:888]),
    .in0(in_reg_wire_2[47]),
    .in1(in_reg_wire_2[111]),
    .in2(in_reg_wire_2[175]),
    .in3(in_reg_wire_2[239]),
    .out0(in_reg_wire_3[188]),
    .out1(in_reg_wire_3[189]),
    .out2(in_reg_wire_3[190]),
    .out3(in_reg_wire_3[191])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_48
  (
    .sel(conf_out[903:896]),
    .in0(in_reg_wire_2[48]),
    .in1(in_reg_wire_2[112]),
    .in2(in_reg_wire_2[176]),
    .in3(in_reg_wire_2[240]),
    .out0(in_reg_wire_3[192]),
    .out1(in_reg_wire_3[193]),
    .out2(in_reg_wire_3[194]),
    .out3(in_reg_wire_3[195])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_49
  (
    .sel(conf_out[911:904]),
    .in0(in_reg_wire_2[49]),
    .in1(in_reg_wire_2[113]),
    .in2(in_reg_wire_2[177]),
    .in3(in_reg_wire_2[241]),
    .out0(in_reg_wire_3[196]),
    .out1(in_reg_wire_3[197]),
    .out2(in_reg_wire_3[198]),
    .out3(in_reg_wire_3[199])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_50
  (
    .sel(conf_out[919:912]),
    .in0(in_reg_wire_2[50]),
    .in1(in_reg_wire_2[114]),
    .in2(in_reg_wire_2[178]),
    .in3(in_reg_wire_2[242]),
    .out0(in_reg_wire_3[200]),
    .out1(in_reg_wire_3[201]),
    .out2(in_reg_wire_3[202]),
    .out3(in_reg_wire_3[203])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_51
  (
    .sel(conf_out[927:920]),
    .in0(in_reg_wire_2[51]),
    .in1(in_reg_wire_2[115]),
    .in2(in_reg_wire_2[179]),
    .in3(in_reg_wire_2[243]),
    .out0(in_reg_wire_3[204]),
    .out1(in_reg_wire_3[205]),
    .out2(in_reg_wire_3[206]),
    .out3(in_reg_wire_3[207])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_52
  (
    .sel(conf_out[935:928]),
    .in0(in_reg_wire_2[52]),
    .in1(in_reg_wire_2[116]),
    .in2(in_reg_wire_2[180]),
    .in3(in_reg_wire_2[244]),
    .out0(in_reg_wire_3[208]),
    .out1(in_reg_wire_3[209]),
    .out2(in_reg_wire_3[210]),
    .out3(in_reg_wire_3[211])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_53
  (
    .sel(conf_out[943:936]),
    .in0(in_reg_wire_2[53]),
    .in1(in_reg_wire_2[117]),
    .in2(in_reg_wire_2[181]),
    .in3(in_reg_wire_2[245]),
    .out0(in_reg_wire_3[212]),
    .out1(in_reg_wire_3[213]),
    .out2(in_reg_wire_3[214]),
    .out3(in_reg_wire_3[215])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_54
  (
    .sel(conf_out[951:944]),
    .in0(in_reg_wire_2[54]),
    .in1(in_reg_wire_2[118]),
    .in2(in_reg_wire_2[182]),
    .in3(in_reg_wire_2[246]),
    .out0(in_reg_wire_3[216]),
    .out1(in_reg_wire_3[217]),
    .out2(in_reg_wire_3[218]),
    .out3(in_reg_wire_3[219])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_55
  (
    .sel(conf_out[959:952]),
    .in0(in_reg_wire_2[55]),
    .in1(in_reg_wire_2[119]),
    .in2(in_reg_wire_2[183]),
    .in3(in_reg_wire_2[247]),
    .out0(in_reg_wire_3[220]),
    .out1(in_reg_wire_3[221]),
    .out2(in_reg_wire_3[222]),
    .out3(in_reg_wire_3[223])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_56
  (
    .sel(conf_out[967:960]),
    .in0(in_reg_wire_2[56]),
    .in1(in_reg_wire_2[120]),
    .in2(in_reg_wire_2[184]),
    .in3(in_reg_wire_2[248]),
    .out0(in_reg_wire_3[224]),
    .out1(in_reg_wire_3[225]),
    .out2(in_reg_wire_3[226]),
    .out3(in_reg_wire_3[227])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_57
  (
    .sel(conf_out[975:968]),
    .in0(in_reg_wire_2[57]),
    .in1(in_reg_wire_2[121]),
    .in2(in_reg_wire_2[185]),
    .in3(in_reg_wire_2[249]),
    .out0(in_reg_wire_3[228]),
    .out1(in_reg_wire_3[229]),
    .out2(in_reg_wire_3[230]),
    .out3(in_reg_wire_3[231])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_58
  (
    .sel(conf_out[983:976]),
    .in0(in_reg_wire_2[58]),
    .in1(in_reg_wire_2[122]),
    .in2(in_reg_wire_2[186]),
    .in3(in_reg_wire_2[250]),
    .out0(in_reg_wire_3[232]),
    .out1(in_reg_wire_3[233]),
    .out2(in_reg_wire_3[234]),
    .out3(in_reg_wire_3[235])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_59
  (
    .sel(conf_out[991:984]),
    .in0(in_reg_wire_2[59]),
    .in1(in_reg_wire_2[123]),
    .in2(in_reg_wire_2[187]),
    .in3(in_reg_wire_2[251]),
    .out0(in_reg_wire_3[236]),
    .out1(in_reg_wire_3[237]),
    .out2(in_reg_wire_3[238]),
    .out3(in_reg_wire_3[239])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_60
  (
    .sel(conf_out[999:992]),
    .in0(in_reg_wire_2[60]),
    .in1(in_reg_wire_2[124]),
    .in2(in_reg_wire_2[188]),
    .in3(in_reg_wire_2[252]),
    .out0(in_reg_wire_3[240]),
    .out1(in_reg_wire_3[241]),
    .out2(in_reg_wire_3[242]),
    .out3(in_reg_wire_3[243])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_61
  (
    .sel(conf_out[1007:1000]),
    .in0(in_reg_wire_2[61]),
    .in1(in_reg_wire_2[125]),
    .in2(in_reg_wire_2[189]),
    .in3(in_reg_wire_2[253]),
    .out0(in_reg_wire_3[244]),
    .out1(in_reg_wire_3[245]),
    .out2(in_reg_wire_3[246]),
    .out3(in_reg_wire_3[247])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_62
  (
    .sel(conf_out[1015:1008]),
    .in0(in_reg_wire_2[62]),
    .in1(in_reg_wire_2[126]),
    .in2(in_reg_wire_2[190]),
    .in3(in_reg_wire_2[254]),
    .out0(in_reg_wire_3[248]),
    .out1(in_reg_wire_3[249]),
    .out2(in_reg_wire_3[250]),
    .out3(in_reg_wire_3[251])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_1_63
  (
    .sel(conf_out[1023:1016]),
    .in0(in_reg_wire_2[63]),
    .in1(in_reg_wire_2[127]),
    .in2(in_reg_wire_2[191]),
    .in3(in_reg_wire_2[255]),
    .out0(in_reg_wire_3[252]),
    .out1(in_reg_wire_3[253]),
    .out2(in_reg_wire_3[254]),
    .out3(in_reg_wire_3[255])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_0
  (
    .sel(conf_out[1031:1024]),
    .in0(in_reg_wire_4[0]),
    .in1(in_reg_wire_4[64]),
    .in2(in_reg_wire_4[128]),
    .in3(in_reg_wire_4[192]),
    .out0(in_reg_wire_5[0]),
    .out1(in_reg_wire_5[1]),
    .out2(in_reg_wire_5[2]),
    .out3(in_reg_wire_5[3])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_1
  (
    .sel(conf_out[1039:1032]),
    .in0(in_reg_wire_4[1]),
    .in1(in_reg_wire_4[65]),
    .in2(in_reg_wire_4[129]),
    .in3(in_reg_wire_4[193]),
    .out0(in_reg_wire_5[4]),
    .out1(in_reg_wire_5[5]),
    .out2(in_reg_wire_5[6]),
    .out3(in_reg_wire_5[7])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_2
  (
    .sel(conf_out[1047:1040]),
    .in0(in_reg_wire_4[2]),
    .in1(in_reg_wire_4[66]),
    .in2(in_reg_wire_4[130]),
    .in3(in_reg_wire_4[194]),
    .out0(in_reg_wire_5[8]),
    .out1(in_reg_wire_5[9]),
    .out2(in_reg_wire_5[10]),
    .out3(in_reg_wire_5[11])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_3
  (
    .sel(conf_out[1055:1048]),
    .in0(in_reg_wire_4[3]),
    .in1(in_reg_wire_4[67]),
    .in2(in_reg_wire_4[131]),
    .in3(in_reg_wire_4[195]),
    .out0(in_reg_wire_5[12]),
    .out1(in_reg_wire_5[13]),
    .out2(in_reg_wire_5[14]),
    .out3(in_reg_wire_5[15])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_4
  (
    .sel(conf_out[1063:1056]),
    .in0(in_reg_wire_4[4]),
    .in1(in_reg_wire_4[68]),
    .in2(in_reg_wire_4[132]),
    .in3(in_reg_wire_4[196]),
    .out0(in_reg_wire_5[16]),
    .out1(in_reg_wire_5[17]),
    .out2(in_reg_wire_5[18]),
    .out3(in_reg_wire_5[19])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_5
  (
    .sel(conf_out[1071:1064]),
    .in0(in_reg_wire_4[5]),
    .in1(in_reg_wire_4[69]),
    .in2(in_reg_wire_4[133]),
    .in3(in_reg_wire_4[197]),
    .out0(in_reg_wire_5[20]),
    .out1(in_reg_wire_5[21]),
    .out2(in_reg_wire_5[22]),
    .out3(in_reg_wire_5[23])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_6
  (
    .sel(conf_out[1079:1072]),
    .in0(in_reg_wire_4[6]),
    .in1(in_reg_wire_4[70]),
    .in2(in_reg_wire_4[134]),
    .in3(in_reg_wire_4[198]),
    .out0(in_reg_wire_5[24]),
    .out1(in_reg_wire_5[25]),
    .out2(in_reg_wire_5[26]),
    .out3(in_reg_wire_5[27])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_7
  (
    .sel(conf_out[1087:1080]),
    .in0(in_reg_wire_4[7]),
    .in1(in_reg_wire_4[71]),
    .in2(in_reg_wire_4[135]),
    .in3(in_reg_wire_4[199]),
    .out0(in_reg_wire_5[28]),
    .out1(in_reg_wire_5[29]),
    .out2(in_reg_wire_5[30]),
    .out3(in_reg_wire_5[31])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_8
  (
    .sel(conf_out[1095:1088]),
    .in0(in_reg_wire_4[8]),
    .in1(in_reg_wire_4[72]),
    .in2(in_reg_wire_4[136]),
    .in3(in_reg_wire_4[200]),
    .out0(in_reg_wire_5[32]),
    .out1(in_reg_wire_5[33]),
    .out2(in_reg_wire_5[34]),
    .out3(in_reg_wire_5[35])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_9
  (
    .sel(conf_out[1103:1096]),
    .in0(in_reg_wire_4[9]),
    .in1(in_reg_wire_4[73]),
    .in2(in_reg_wire_4[137]),
    .in3(in_reg_wire_4[201]),
    .out0(in_reg_wire_5[36]),
    .out1(in_reg_wire_5[37]),
    .out2(in_reg_wire_5[38]),
    .out3(in_reg_wire_5[39])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_10
  (
    .sel(conf_out[1111:1104]),
    .in0(in_reg_wire_4[10]),
    .in1(in_reg_wire_4[74]),
    .in2(in_reg_wire_4[138]),
    .in3(in_reg_wire_4[202]),
    .out0(in_reg_wire_5[40]),
    .out1(in_reg_wire_5[41]),
    .out2(in_reg_wire_5[42]),
    .out3(in_reg_wire_5[43])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_11
  (
    .sel(conf_out[1119:1112]),
    .in0(in_reg_wire_4[11]),
    .in1(in_reg_wire_4[75]),
    .in2(in_reg_wire_4[139]),
    .in3(in_reg_wire_4[203]),
    .out0(in_reg_wire_5[44]),
    .out1(in_reg_wire_5[45]),
    .out2(in_reg_wire_5[46]),
    .out3(in_reg_wire_5[47])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_12
  (
    .sel(conf_out[1127:1120]),
    .in0(in_reg_wire_4[12]),
    .in1(in_reg_wire_4[76]),
    .in2(in_reg_wire_4[140]),
    .in3(in_reg_wire_4[204]),
    .out0(in_reg_wire_5[48]),
    .out1(in_reg_wire_5[49]),
    .out2(in_reg_wire_5[50]),
    .out3(in_reg_wire_5[51])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_13
  (
    .sel(conf_out[1135:1128]),
    .in0(in_reg_wire_4[13]),
    .in1(in_reg_wire_4[77]),
    .in2(in_reg_wire_4[141]),
    .in3(in_reg_wire_4[205]),
    .out0(in_reg_wire_5[52]),
    .out1(in_reg_wire_5[53]),
    .out2(in_reg_wire_5[54]),
    .out3(in_reg_wire_5[55])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_14
  (
    .sel(conf_out[1143:1136]),
    .in0(in_reg_wire_4[14]),
    .in1(in_reg_wire_4[78]),
    .in2(in_reg_wire_4[142]),
    .in3(in_reg_wire_4[206]),
    .out0(in_reg_wire_5[56]),
    .out1(in_reg_wire_5[57]),
    .out2(in_reg_wire_5[58]),
    .out3(in_reg_wire_5[59])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_15
  (
    .sel(conf_out[1151:1144]),
    .in0(in_reg_wire_4[15]),
    .in1(in_reg_wire_4[79]),
    .in2(in_reg_wire_4[143]),
    .in3(in_reg_wire_4[207]),
    .out0(in_reg_wire_5[60]),
    .out1(in_reg_wire_5[61]),
    .out2(in_reg_wire_5[62]),
    .out3(in_reg_wire_5[63])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_16
  (
    .sel(conf_out[1159:1152]),
    .in0(in_reg_wire_4[16]),
    .in1(in_reg_wire_4[80]),
    .in2(in_reg_wire_4[144]),
    .in3(in_reg_wire_4[208]),
    .out0(in_reg_wire_5[64]),
    .out1(in_reg_wire_5[65]),
    .out2(in_reg_wire_5[66]),
    .out3(in_reg_wire_5[67])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_17
  (
    .sel(conf_out[1167:1160]),
    .in0(in_reg_wire_4[17]),
    .in1(in_reg_wire_4[81]),
    .in2(in_reg_wire_4[145]),
    .in3(in_reg_wire_4[209]),
    .out0(in_reg_wire_5[68]),
    .out1(in_reg_wire_5[69]),
    .out2(in_reg_wire_5[70]),
    .out3(in_reg_wire_5[71])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_18
  (
    .sel(conf_out[1175:1168]),
    .in0(in_reg_wire_4[18]),
    .in1(in_reg_wire_4[82]),
    .in2(in_reg_wire_4[146]),
    .in3(in_reg_wire_4[210]),
    .out0(in_reg_wire_5[72]),
    .out1(in_reg_wire_5[73]),
    .out2(in_reg_wire_5[74]),
    .out3(in_reg_wire_5[75])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_19
  (
    .sel(conf_out[1183:1176]),
    .in0(in_reg_wire_4[19]),
    .in1(in_reg_wire_4[83]),
    .in2(in_reg_wire_4[147]),
    .in3(in_reg_wire_4[211]),
    .out0(in_reg_wire_5[76]),
    .out1(in_reg_wire_5[77]),
    .out2(in_reg_wire_5[78]),
    .out3(in_reg_wire_5[79])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_20
  (
    .sel(conf_out[1191:1184]),
    .in0(in_reg_wire_4[20]),
    .in1(in_reg_wire_4[84]),
    .in2(in_reg_wire_4[148]),
    .in3(in_reg_wire_4[212]),
    .out0(in_reg_wire_5[80]),
    .out1(in_reg_wire_5[81]),
    .out2(in_reg_wire_5[82]),
    .out3(in_reg_wire_5[83])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_21
  (
    .sel(conf_out[1199:1192]),
    .in0(in_reg_wire_4[21]),
    .in1(in_reg_wire_4[85]),
    .in2(in_reg_wire_4[149]),
    .in3(in_reg_wire_4[213]),
    .out0(in_reg_wire_5[84]),
    .out1(in_reg_wire_5[85]),
    .out2(in_reg_wire_5[86]),
    .out3(in_reg_wire_5[87])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_22
  (
    .sel(conf_out[1207:1200]),
    .in0(in_reg_wire_4[22]),
    .in1(in_reg_wire_4[86]),
    .in2(in_reg_wire_4[150]),
    .in3(in_reg_wire_4[214]),
    .out0(in_reg_wire_5[88]),
    .out1(in_reg_wire_5[89]),
    .out2(in_reg_wire_5[90]),
    .out3(in_reg_wire_5[91])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_23
  (
    .sel(conf_out[1215:1208]),
    .in0(in_reg_wire_4[23]),
    .in1(in_reg_wire_4[87]),
    .in2(in_reg_wire_4[151]),
    .in3(in_reg_wire_4[215]),
    .out0(in_reg_wire_5[92]),
    .out1(in_reg_wire_5[93]),
    .out2(in_reg_wire_5[94]),
    .out3(in_reg_wire_5[95])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_24
  (
    .sel(conf_out[1223:1216]),
    .in0(in_reg_wire_4[24]),
    .in1(in_reg_wire_4[88]),
    .in2(in_reg_wire_4[152]),
    .in3(in_reg_wire_4[216]),
    .out0(in_reg_wire_5[96]),
    .out1(in_reg_wire_5[97]),
    .out2(in_reg_wire_5[98]),
    .out3(in_reg_wire_5[99])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_25
  (
    .sel(conf_out[1231:1224]),
    .in0(in_reg_wire_4[25]),
    .in1(in_reg_wire_4[89]),
    .in2(in_reg_wire_4[153]),
    .in3(in_reg_wire_4[217]),
    .out0(in_reg_wire_5[100]),
    .out1(in_reg_wire_5[101]),
    .out2(in_reg_wire_5[102]),
    .out3(in_reg_wire_5[103])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_26
  (
    .sel(conf_out[1239:1232]),
    .in0(in_reg_wire_4[26]),
    .in1(in_reg_wire_4[90]),
    .in2(in_reg_wire_4[154]),
    .in3(in_reg_wire_4[218]),
    .out0(in_reg_wire_5[104]),
    .out1(in_reg_wire_5[105]),
    .out2(in_reg_wire_5[106]),
    .out3(in_reg_wire_5[107])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_27
  (
    .sel(conf_out[1247:1240]),
    .in0(in_reg_wire_4[27]),
    .in1(in_reg_wire_4[91]),
    .in2(in_reg_wire_4[155]),
    .in3(in_reg_wire_4[219]),
    .out0(in_reg_wire_5[108]),
    .out1(in_reg_wire_5[109]),
    .out2(in_reg_wire_5[110]),
    .out3(in_reg_wire_5[111])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_28
  (
    .sel(conf_out[1255:1248]),
    .in0(in_reg_wire_4[28]),
    .in1(in_reg_wire_4[92]),
    .in2(in_reg_wire_4[156]),
    .in3(in_reg_wire_4[220]),
    .out0(in_reg_wire_5[112]),
    .out1(in_reg_wire_5[113]),
    .out2(in_reg_wire_5[114]),
    .out3(in_reg_wire_5[115])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_29
  (
    .sel(conf_out[1263:1256]),
    .in0(in_reg_wire_4[29]),
    .in1(in_reg_wire_4[93]),
    .in2(in_reg_wire_4[157]),
    .in3(in_reg_wire_4[221]),
    .out0(in_reg_wire_5[116]),
    .out1(in_reg_wire_5[117]),
    .out2(in_reg_wire_5[118]),
    .out3(in_reg_wire_5[119])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_30
  (
    .sel(conf_out[1271:1264]),
    .in0(in_reg_wire_4[30]),
    .in1(in_reg_wire_4[94]),
    .in2(in_reg_wire_4[158]),
    .in3(in_reg_wire_4[222]),
    .out0(in_reg_wire_5[120]),
    .out1(in_reg_wire_5[121]),
    .out2(in_reg_wire_5[122]),
    .out3(in_reg_wire_5[123])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_31
  (
    .sel(conf_out[1279:1272]),
    .in0(in_reg_wire_4[31]),
    .in1(in_reg_wire_4[95]),
    .in2(in_reg_wire_4[159]),
    .in3(in_reg_wire_4[223]),
    .out0(in_reg_wire_5[124]),
    .out1(in_reg_wire_5[125]),
    .out2(in_reg_wire_5[126]),
    .out3(in_reg_wire_5[127])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_32
  (
    .sel(conf_out[1287:1280]),
    .in0(in_reg_wire_4[32]),
    .in1(in_reg_wire_4[96]),
    .in2(in_reg_wire_4[160]),
    .in3(in_reg_wire_4[224]),
    .out0(in_reg_wire_5[128]),
    .out1(in_reg_wire_5[129]),
    .out2(in_reg_wire_5[130]),
    .out3(in_reg_wire_5[131])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_33
  (
    .sel(conf_out[1295:1288]),
    .in0(in_reg_wire_4[33]),
    .in1(in_reg_wire_4[97]),
    .in2(in_reg_wire_4[161]),
    .in3(in_reg_wire_4[225]),
    .out0(in_reg_wire_5[132]),
    .out1(in_reg_wire_5[133]),
    .out2(in_reg_wire_5[134]),
    .out3(in_reg_wire_5[135])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_34
  (
    .sel(conf_out[1303:1296]),
    .in0(in_reg_wire_4[34]),
    .in1(in_reg_wire_4[98]),
    .in2(in_reg_wire_4[162]),
    .in3(in_reg_wire_4[226]),
    .out0(in_reg_wire_5[136]),
    .out1(in_reg_wire_5[137]),
    .out2(in_reg_wire_5[138]),
    .out3(in_reg_wire_5[139])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_35
  (
    .sel(conf_out[1311:1304]),
    .in0(in_reg_wire_4[35]),
    .in1(in_reg_wire_4[99]),
    .in2(in_reg_wire_4[163]),
    .in3(in_reg_wire_4[227]),
    .out0(in_reg_wire_5[140]),
    .out1(in_reg_wire_5[141]),
    .out2(in_reg_wire_5[142]),
    .out3(in_reg_wire_5[143])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_36
  (
    .sel(conf_out[1319:1312]),
    .in0(in_reg_wire_4[36]),
    .in1(in_reg_wire_4[100]),
    .in2(in_reg_wire_4[164]),
    .in3(in_reg_wire_4[228]),
    .out0(in_reg_wire_5[144]),
    .out1(in_reg_wire_5[145]),
    .out2(in_reg_wire_5[146]),
    .out3(in_reg_wire_5[147])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_37
  (
    .sel(conf_out[1327:1320]),
    .in0(in_reg_wire_4[37]),
    .in1(in_reg_wire_4[101]),
    .in2(in_reg_wire_4[165]),
    .in3(in_reg_wire_4[229]),
    .out0(in_reg_wire_5[148]),
    .out1(in_reg_wire_5[149]),
    .out2(in_reg_wire_5[150]),
    .out3(in_reg_wire_5[151])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_38
  (
    .sel(conf_out[1335:1328]),
    .in0(in_reg_wire_4[38]),
    .in1(in_reg_wire_4[102]),
    .in2(in_reg_wire_4[166]),
    .in3(in_reg_wire_4[230]),
    .out0(in_reg_wire_5[152]),
    .out1(in_reg_wire_5[153]),
    .out2(in_reg_wire_5[154]),
    .out3(in_reg_wire_5[155])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_39
  (
    .sel(conf_out[1343:1336]),
    .in0(in_reg_wire_4[39]),
    .in1(in_reg_wire_4[103]),
    .in2(in_reg_wire_4[167]),
    .in3(in_reg_wire_4[231]),
    .out0(in_reg_wire_5[156]),
    .out1(in_reg_wire_5[157]),
    .out2(in_reg_wire_5[158]),
    .out3(in_reg_wire_5[159])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_40
  (
    .sel(conf_out[1351:1344]),
    .in0(in_reg_wire_4[40]),
    .in1(in_reg_wire_4[104]),
    .in2(in_reg_wire_4[168]),
    .in3(in_reg_wire_4[232]),
    .out0(in_reg_wire_5[160]),
    .out1(in_reg_wire_5[161]),
    .out2(in_reg_wire_5[162]),
    .out3(in_reg_wire_5[163])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_41
  (
    .sel(conf_out[1359:1352]),
    .in0(in_reg_wire_4[41]),
    .in1(in_reg_wire_4[105]),
    .in2(in_reg_wire_4[169]),
    .in3(in_reg_wire_4[233]),
    .out0(in_reg_wire_5[164]),
    .out1(in_reg_wire_5[165]),
    .out2(in_reg_wire_5[166]),
    .out3(in_reg_wire_5[167])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_42
  (
    .sel(conf_out[1367:1360]),
    .in0(in_reg_wire_4[42]),
    .in1(in_reg_wire_4[106]),
    .in2(in_reg_wire_4[170]),
    .in3(in_reg_wire_4[234]),
    .out0(in_reg_wire_5[168]),
    .out1(in_reg_wire_5[169]),
    .out2(in_reg_wire_5[170]),
    .out3(in_reg_wire_5[171])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_43
  (
    .sel(conf_out[1375:1368]),
    .in0(in_reg_wire_4[43]),
    .in1(in_reg_wire_4[107]),
    .in2(in_reg_wire_4[171]),
    .in3(in_reg_wire_4[235]),
    .out0(in_reg_wire_5[172]),
    .out1(in_reg_wire_5[173]),
    .out2(in_reg_wire_5[174]),
    .out3(in_reg_wire_5[175])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_44
  (
    .sel(conf_out[1383:1376]),
    .in0(in_reg_wire_4[44]),
    .in1(in_reg_wire_4[108]),
    .in2(in_reg_wire_4[172]),
    .in3(in_reg_wire_4[236]),
    .out0(in_reg_wire_5[176]),
    .out1(in_reg_wire_5[177]),
    .out2(in_reg_wire_5[178]),
    .out3(in_reg_wire_5[179])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_45
  (
    .sel(conf_out[1391:1384]),
    .in0(in_reg_wire_4[45]),
    .in1(in_reg_wire_4[109]),
    .in2(in_reg_wire_4[173]),
    .in3(in_reg_wire_4[237]),
    .out0(in_reg_wire_5[180]),
    .out1(in_reg_wire_5[181]),
    .out2(in_reg_wire_5[182]),
    .out3(in_reg_wire_5[183])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_46
  (
    .sel(conf_out[1399:1392]),
    .in0(in_reg_wire_4[46]),
    .in1(in_reg_wire_4[110]),
    .in2(in_reg_wire_4[174]),
    .in3(in_reg_wire_4[238]),
    .out0(in_reg_wire_5[184]),
    .out1(in_reg_wire_5[185]),
    .out2(in_reg_wire_5[186]),
    .out3(in_reg_wire_5[187])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_47
  (
    .sel(conf_out[1407:1400]),
    .in0(in_reg_wire_4[47]),
    .in1(in_reg_wire_4[111]),
    .in2(in_reg_wire_4[175]),
    .in3(in_reg_wire_4[239]),
    .out0(in_reg_wire_5[188]),
    .out1(in_reg_wire_5[189]),
    .out2(in_reg_wire_5[190]),
    .out3(in_reg_wire_5[191])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_48
  (
    .sel(conf_out[1415:1408]),
    .in0(in_reg_wire_4[48]),
    .in1(in_reg_wire_4[112]),
    .in2(in_reg_wire_4[176]),
    .in3(in_reg_wire_4[240]),
    .out0(in_reg_wire_5[192]),
    .out1(in_reg_wire_5[193]),
    .out2(in_reg_wire_5[194]),
    .out3(in_reg_wire_5[195])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_49
  (
    .sel(conf_out[1423:1416]),
    .in0(in_reg_wire_4[49]),
    .in1(in_reg_wire_4[113]),
    .in2(in_reg_wire_4[177]),
    .in3(in_reg_wire_4[241]),
    .out0(in_reg_wire_5[196]),
    .out1(in_reg_wire_5[197]),
    .out2(in_reg_wire_5[198]),
    .out3(in_reg_wire_5[199])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_50
  (
    .sel(conf_out[1431:1424]),
    .in0(in_reg_wire_4[50]),
    .in1(in_reg_wire_4[114]),
    .in2(in_reg_wire_4[178]),
    .in3(in_reg_wire_4[242]),
    .out0(in_reg_wire_5[200]),
    .out1(in_reg_wire_5[201]),
    .out2(in_reg_wire_5[202]),
    .out3(in_reg_wire_5[203])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_51
  (
    .sel(conf_out[1439:1432]),
    .in0(in_reg_wire_4[51]),
    .in1(in_reg_wire_4[115]),
    .in2(in_reg_wire_4[179]),
    .in3(in_reg_wire_4[243]),
    .out0(in_reg_wire_5[204]),
    .out1(in_reg_wire_5[205]),
    .out2(in_reg_wire_5[206]),
    .out3(in_reg_wire_5[207])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_52
  (
    .sel(conf_out[1447:1440]),
    .in0(in_reg_wire_4[52]),
    .in1(in_reg_wire_4[116]),
    .in2(in_reg_wire_4[180]),
    .in3(in_reg_wire_4[244]),
    .out0(in_reg_wire_5[208]),
    .out1(in_reg_wire_5[209]),
    .out2(in_reg_wire_5[210]),
    .out3(in_reg_wire_5[211])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_53
  (
    .sel(conf_out[1455:1448]),
    .in0(in_reg_wire_4[53]),
    .in1(in_reg_wire_4[117]),
    .in2(in_reg_wire_4[181]),
    .in3(in_reg_wire_4[245]),
    .out0(in_reg_wire_5[212]),
    .out1(in_reg_wire_5[213]),
    .out2(in_reg_wire_5[214]),
    .out3(in_reg_wire_5[215])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_54
  (
    .sel(conf_out[1463:1456]),
    .in0(in_reg_wire_4[54]),
    .in1(in_reg_wire_4[118]),
    .in2(in_reg_wire_4[182]),
    .in3(in_reg_wire_4[246]),
    .out0(in_reg_wire_5[216]),
    .out1(in_reg_wire_5[217]),
    .out2(in_reg_wire_5[218]),
    .out3(in_reg_wire_5[219])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_55
  (
    .sel(conf_out[1471:1464]),
    .in0(in_reg_wire_4[55]),
    .in1(in_reg_wire_4[119]),
    .in2(in_reg_wire_4[183]),
    .in3(in_reg_wire_4[247]),
    .out0(in_reg_wire_5[220]),
    .out1(in_reg_wire_5[221]),
    .out2(in_reg_wire_5[222]),
    .out3(in_reg_wire_5[223])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_56
  (
    .sel(conf_out[1479:1472]),
    .in0(in_reg_wire_4[56]),
    .in1(in_reg_wire_4[120]),
    .in2(in_reg_wire_4[184]),
    .in3(in_reg_wire_4[248]),
    .out0(in_reg_wire_5[224]),
    .out1(in_reg_wire_5[225]),
    .out2(in_reg_wire_5[226]),
    .out3(in_reg_wire_5[227])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_57
  (
    .sel(conf_out[1487:1480]),
    .in0(in_reg_wire_4[57]),
    .in1(in_reg_wire_4[121]),
    .in2(in_reg_wire_4[185]),
    .in3(in_reg_wire_4[249]),
    .out0(in_reg_wire_5[228]),
    .out1(in_reg_wire_5[229]),
    .out2(in_reg_wire_5[230]),
    .out3(in_reg_wire_5[231])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_58
  (
    .sel(conf_out[1495:1488]),
    .in0(in_reg_wire_4[58]),
    .in1(in_reg_wire_4[122]),
    .in2(in_reg_wire_4[186]),
    .in3(in_reg_wire_4[250]),
    .out0(in_reg_wire_5[232]),
    .out1(in_reg_wire_5[233]),
    .out2(in_reg_wire_5[234]),
    .out3(in_reg_wire_5[235])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_59
  (
    .sel(conf_out[1503:1496]),
    .in0(in_reg_wire_4[59]),
    .in1(in_reg_wire_4[123]),
    .in2(in_reg_wire_4[187]),
    .in3(in_reg_wire_4[251]),
    .out0(in_reg_wire_5[236]),
    .out1(in_reg_wire_5[237]),
    .out2(in_reg_wire_5[238]),
    .out3(in_reg_wire_5[239])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_60
  (
    .sel(conf_out[1511:1504]),
    .in0(in_reg_wire_4[60]),
    .in1(in_reg_wire_4[124]),
    .in2(in_reg_wire_4[188]),
    .in3(in_reg_wire_4[252]),
    .out0(in_reg_wire_5[240]),
    .out1(in_reg_wire_5[241]),
    .out2(in_reg_wire_5[242]),
    .out3(in_reg_wire_5[243])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_61
  (
    .sel(conf_out[1519:1512]),
    .in0(in_reg_wire_4[61]),
    .in1(in_reg_wire_4[125]),
    .in2(in_reg_wire_4[189]),
    .in3(in_reg_wire_4[253]),
    .out0(in_reg_wire_5[244]),
    .out1(in_reg_wire_5[245]),
    .out2(in_reg_wire_5[246]),
    .out3(in_reg_wire_5[247])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_62
  (
    .sel(conf_out[1527:1520]),
    .in0(in_reg_wire_4[62]),
    .in1(in_reg_wire_4[126]),
    .in2(in_reg_wire_4[190]),
    .in3(in_reg_wire_4[254]),
    .out0(in_reg_wire_5[248]),
    .out1(in_reg_wire_5[249]),
    .out2(in_reg_wire_5[250]),
    .out3(in_reg_wire_5[251])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_2_63
  (
    .sel(conf_out[1535:1528]),
    .in0(in_reg_wire_4[63]),
    .in1(in_reg_wire_4[127]),
    .in2(in_reg_wire_4[191]),
    .in3(in_reg_wire_4[255]),
    .out0(in_reg_wire_5[252]),
    .out1(in_reg_wire_5[253]),
    .out2(in_reg_wire_5[254]),
    .out3(in_reg_wire_5[255])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_0
  (
    .sel(conf_out[1543:1536]),
    .in0(in_reg_wire_6[0]),
    .in1(in_reg_wire_6[64]),
    .in2(in_reg_wire_6[128]),
    .in3(in_reg_wire_6[192]),
    .out0(in_reg_wire_7[0]),
    .out1(in_reg_wire_7[1]),
    .out2(in_reg_wire_7[2]),
    .out3(in_reg_wire_7[3])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_1
  (
    .sel(conf_out[1551:1544]),
    .in0(in_reg_wire_6[1]),
    .in1(in_reg_wire_6[65]),
    .in2(in_reg_wire_6[129]),
    .in3(in_reg_wire_6[193]),
    .out0(in_reg_wire_7[4]),
    .out1(in_reg_wire_7[5]),
    .out2(in_reg_wire_7[6]),
    .out3(in_reg_wire_7[7])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_2
  (
    .sel(conf_out[1559:1552]),
    .in0(in_reg_wire_6[2]),
    .in1(in_reg_wire_6[66]),
    .in2(in_reg_wire_6[130]),
    .in3(in_reg_wire_6[194]),
    .out0(in_reg_wire_7[8]),
    .out1(in_reg_wire_7[9]),
    .out2(in_reg_wire_7[10]),
    .out3(in_reg_wire_7[11])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_3
  (
    .sel(conf_out[1567:1560]),
    .in0(in_reg_wire_6[3]),
    .in1(in_reg_wire_6[67]),
    .in2(in_reg_wire_6[131]),
    .in3(in_reg_wire_6[195]),
    .out0(in_reg_wire_7[12]),
    .out1(in_reg_wire_7[13]),
    .out2(in_reg_wire_7[14]),
    .out3(in_reg_wire_7[15])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_4
  (
    .sel(conf_out[1575:1568]),
    .in0(in_reg_wire_6[4]),
    .in1(in_reg_wire_6[68]),
    .in2(in_reg_wire_6[132]),
    .in3(in_reg_wire_6[196]),
    .out0(in_reg_wire_7[16]),
    .out1(in_reg_wire_7[17]),
    .out2(in_reg_wire_7[18]),
    .out3(in_reg_wire_7[19])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_5
  (
    .sel(conf_out[1583:1576]),
    .in0(in_reg_wire_6[5]),
    .in1(in_reg_wire_6[69]),
    .in2(in_reg_wire_6[133]),
    .in3(in_reg_wire_6[197]),
    .out0(in_reg_wire_7[20]),
    .out1(in_reg_wire_7[21]),
    .out2(in_reg_wire_7[22]),
    .out3(in_reg_wire_7[23])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_6
  (
    .sel(conf_out[1591:1584]),
    .in0(in_reg_wire_6[6]),
    .in1(in_reg_wire_6[70]),
    .in2(in_reg_wire_6[134]),
    .in3(in_reg_wire_6[198]),
    .out0(in_reg_wire_7[24]),
    .out1(in_reg_wire_7[25]),
    .out2(in_reg_wire_7[26]),
    .out3(in_reg_wire_7[27])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_7
  (
    .sel(conf_out[1599:1592]),
    .in0(in_reg_wire_6[7]),
    .in1(in_reg_wire_6[71]),
    .in2(in_reg_wire_6[135]),
    .in3(in_reg_wire_6[199]),
    .out0(in_reg_wire_7[28]),
    .out1(in_reg_wire_7[29]),
    .out2(in_reg_wire_7[30]),
    .out3(in_reg_wire_7[31])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_8
  (
    .sel(conf_out[1607:1600]),
    .in0(in_reg_wire_6[8]),
    .in1(in_reg_wire_6[72]),
    .in2(in_reg_wire_6[136]),
    .in3(in_reg_wire_6[200]),
    .out0(in_reg_wire_7[32]),
    .out1(in_reg_wire_7[33]),
    .out2(in_reg_wire_7[34]),
    .out3(in_reg_wire_7[35])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_9
  (
    .sel(conf_out[1615:1608]),
    .in0(in_reg_wire_6[9]),
    .in1(in_reg_wire_6[73]),
    .in2(in_reg_wire_6[137]),
    .in3(in_reg_wire_6[201]),
    .out0(in_reg_wire_7[36]),
    .out1(in_reg_wire_7[37]),
    .out2(in_reg_wire_7[38]),
    .out3(in_reg_wire_7[39])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_10
  (
    .sel(conf_out[1623:1616]),
    .in0(in_reg_wire_6[10]),
    .in1(in_reg_wire_6[74]),
    .in2(in_reg_wire_6[138]),
    .in3(in_reg_wire_6[202]),
    .out0(in_reg_wire_7[40]),
    .out1(in_reg_wire_7[41]),
    .out2(in_reg_wire_7[42]),
    .out3(in_reg_wire_7[43])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_11
  (
    .sel(conf_out[1631:1624]),
    .in0(in_reg_wire_6[11]),
    .in1(in_reg_wire_6[75]),
    .in2(in_reg_wire_6[139]),
    .in3(in_reg_wire_6[203]),
    .out0(in_reg_wire_7[44]),
    .out1(in_reg_wire_7[45]),
    .out2(in_reg_wire_7[46]),
    .out3(in_reg_wire_7[47])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_12
  (
    .sel(conf_out[1639:1632]),
    .in0(in_reg_wire_6[12]),
    .in1(in_reg_wire_6[76]),
    .in2(in_reg_wire_6[140]),
    .in3(in_reg_wire_6[204]),
    .out0(in_reg_wire_7[48]),
    .out1(in_reg_wire_7[49]),
    .out2(in_reg_wire_7[50]),
    .out3(in_reg_wire_7[51])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_13
  (
    .sel(conf_out[1647:1640]),
    .in0(in_reg_wire_6[13]),
    .in1(in_reg_wire_6[77]),
    .in2(in_reg_wire_6[141]),
    .in3(in_reg_wire_6[205]),
    .out0(in_reg_wire_7[52]),
    .out1(in_reg_wire_7[53]),
    .out2(in_reg_wire_7[54]),
    .out3(in_reg_wire_7[55])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_14
  (
    .sel(conf_out[1655:1648]),
    .in0(in_reg_wire_6[14]),
    .in1(in_reg_wire_6[78]),
    .in2(in_reg_wire_6[142]),
    .in3(in_reg_wire_6[206]),
    .out0(in_reg_wire_7[56]),
    .out1(in_reg_wire_7[57]),
    .out2(in_reg_wire_7[58]),
    .out3(in_reg_wire_7[59])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_15
  (
    .sel(conf_out[1663:1656]),
    .in0(in_reg_wire_6[15]),
    .in1(in_reg_wire_6[79]),
    .in2(in_reg_wire_6[143]),
    .in3(in_reg_wire_6[207]),
    .out0(in_reg_wire_7[60]),
    .out1(in_reg_wire_7[61]),
    .out2(in_reg_wire_7[62]),
    .out3(in_reg_wire_7[63])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_16
  (
    .sel(conf_out[1671:1664]),
    .in0(in_reg_wire_6[16]),
    .in1(in_reg_wire_6[80]),
    .in2(in_reg_wire_6[144]),
    .in3(in_reg_wire_6[208]),
    .out0(in_reg_wire_7[64]),
    .out1(in_reg_wire_7[65]),
    .out2(in_reg_wire_7[66]),
    .out3(in_reg_wire_7[67])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_17
  (
    .sel(conf_out[1679:1672]),
    .in0(in_reg_wire_6[17]),
    .in1(in_reg_wire_6[81]),
    .in2(in_reg_wire_6[145]),
    .in3(in_reg_wire_6[209]),
    .out0(in_reg_wire_7[68]),
    .out1(in_reg_wire_7[69]),
    .out2(in_reg_wire_7[70]),
    .out3(in_reg_wire_7[71])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_18
  (
    .sel(conf_out[1687:1680]),
    .in0(in_reg_wire_6[18]),
    .in1(in_reg_wire_6[82]),
    .in2(in_reg_wire_6[146]),
    .in3(in_reg_wire_6[210]),
    .out0(in_reg_wire_7[72]),
    .out1(in_reg_wire_7[73]),
    .out2(in_reg_wire_7[74]),
    .out3(in_reg_wire_7[75])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_19
  (
    .sel(conf_out[1695:1688]),
    .in0(in_reg_wire_6[19]),
    .in1(in_reg_wire_6[83]),
    .in2(in_reg_wire_6[147]),
    .in3(in_reg_wire_6[211]),
    .out0(in_reg_wire_7[76]),
    .out1(in_reg_wire_7[77]),
    .out2(in_reg_wire_7[78]),
    .out3(in_reg_wire_7[79])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_20
  (
    .sel(conf_out[1703:1696]),
    .in0(in_reg_wire_6[20]),
    .in1(in_reg_wire_6[84]),
    .in2(in_reg_wire_6[148]),
    .in3(in_reg_wire_6[212]),
    .out0(in_reg_wire_7[80]),
    .out1(in_reg_wire_7[81]),
    .out2(in_reg_wire_7[82]),
    .out3(in_reg_wire_7[83])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_21
  (
    .sel(conf_out[1711:1704]),
    .in0(in_reg_wire_6[21]),
    .in1(in_reg_wire_6[85]),
    .in2(in_reg_wire_6[149]),
    .in3(in_reg_wire_6[213]),
    .out0(in_reg_wire_7[84]),
    .out1(in_reg_wire_7[85]),
    .out2(in_reg_wire_7[86]),
    .out3(in_reg_wire_7[87])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_22
  (
    .sel(conf_out[1719:1712]),
    .in0(in_reg_wire_6[22]),
    .in1(in_reg_wire_6[86]),
    .in2(in_reg_wire_6[150]),
    .in3(in_reg_wire_6[214]),
    .out0(in_reg_wire_7[88]),
    .out1(in_reg_wire_7[89]),
    .out2(in_reg_wire_7[90]),
    .out3(in_reg_wire_7[91])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_23
  (
    .sel(conf_out[1727:1720]),
    .in0(in_reg_wire_6[23]),
    .in1(in_reg_wire_6[87]),
    .in2(in_reg_wire_6[151]),
    .in3(in_reg_wire_6[215]),
    .out0(in_reg_wire_7[92]),
    .out1(in_reg_wire_7[93]),
    .out2(in_reg_wire_7[94]),
    .out3(in_reg_wire_7[95])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_24
  (
    .sel(conf_out[1735:1728]),
    .in0(in_reg_wire_6[24]),
    .in1(in_reg_wire_6[88]),
    .in2(in_reg_wire_6[152]),
    .in3(in_reg_wire_6[216]),
    .out0(in_reg_wire_7[96]),
    .out1(in_reg_wire_7[97]),
    .out2(in_reg_wire_7[98]),
    .out3(in_reg_wire_7[99])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_25
  (
    .sel(conf_out[1743:1736]),
    .in0(in_reg_wire_6[25]),
    .in1(in_reg_wire_6[89]),
    .in2(in_reg_wire_6[153]),
    .in3(in_reg_wire_6[217]),
    .out0(in_reg_wire_7[100]),
    .out1(in_reg_wire_7[101]),
    .out2(in_reg_wire_7[102]),
    .out3(in_reg_wire_7[103])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_26
  (
    .sel(conf_out[1751:1744]),
    .in0(in_reg_wire_6[26]),
    .in1(in_reg_wire_6[90]),
    .in2(in_reg_wire_6[154]),
    .in3(in_reg_wire_6[218]),
    .out0(in_reg_wire_7[104]),
    .out1(in_reg_wire_7[105]),
    .out2(in_reg_wire_7[106]),
    .out3(in_reg_wire_7[107])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_27
  (
    .sel(conf_out[1759:1752]),
    .in0(in_reg_wire_6[27]),
    .in1(in_reg_wire_6[91]),
    .in2(in_reg_wire_6[155]),
    .in3(in_reg_wire_6[219]),
    .out0(in_reg_wire_7[108]),
    .out1(in_reg_wire_7[109]),
    .out2(in_reg_wire_7[110]),
    .out3(in_reg_wire_7[111])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_28
  (
    .sel(conf_out[1767:1760]),
    .in0(in_reg_wire_6[28]),
    .in1(in_reg_wire_6[92]),
    .in2(in_reg_wire_6[156]),
    .in3(in_reg_wire_6[220]),
    .out0(in_reg_wire_7[112]),
    .out1(in_reg_wire_7[113]),
    .out2(in_reg_wire_7[114]),
    .out3(in_reg_wire_7[115])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_29
  (
    .sel(conf_out[1775:1768]),
    .in0(in_reg_wire_6[29]),
    .in1(in_reg_wire_6[93]),
    .in2(in_reg_wire_6[157]),
    .in3(in_reg_wire_6[221]),
    .out0(in_reg_wire_7[116]),
    .out1(in_reg_wire_7[117]),
    .out2(in_reg_wire_7[118]),
    .out3(in_reg_wire_7[119])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_30
  (
    .sel(conf_out[1783:1776]),
    .in0(in_reg_wire_6[30]),
    .in1(in_reg_wire_6[94]),
    .in2(in_reg_wire_6[158]),
    .in3(in_reg_wire_6[222]),
    .out0(in_reg_wire_7[120]),
    .out1(in_reg_wire_7[121]),
    .out2(in_reg_wire_7[122]),
    .out3(in_reg_wire_7[123])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_31
  (
    .sel(conf_out[1791:1784]),
    .in0(in_reg_wire_6[31]),
    .in1(in_reg_wire_6[95]),
    .in2(in_reg_wire_6[159]),
    .in3(in_reg_wire_6[223]),
    .out0(in_reg_wire_7[124]),
    .out1(in_reg_wire_7[125]),
    .out2(in_reg_wire_7[126]),
    .out3(in_reg_wire_7[127])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_32
  (
    .sel(conf_out[1799:1792]),
    .in0(in_reg_wire_6[32]),
    .in1(in_reg_wire_6[96]),
    .in2(in_reg_wire_6[160]),
    .in3(in_reg_wire_6[224]),
    .out0(in_reg_wire_7[128]),
    .out1(in_reg_wire_7[129]),
    .out2(in_reg_wire_7[130]),
    .out3(in_reg_wire_7[131])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_33
  (
    .sel(conf_out[1807:1800]),
    .in0(in_reg_wire_6[33]),
    .in1(in_reg_wire_6[97]),
    .in2(in_reg_wire_6[161]),
    .in3(in_reg_wire_6[225]),
    .out0(in_reg_wire_7[132]),
    .out1(in_reg_wire_7[133]),
    .out2(in_reg_wire_7[134]),
    .out3(in_reg_wire_7[135])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_34
  (
    .sel(conf_out[1815:1808]),
    .in0(in_reg_wire_6[34]),
    .in1(in_reg_wire_6[98]),
    .in2(in_reg_wire_6[162]),
    .in3(in_reg_wire_6[226]),
    .out0(in_reg_wire_7[136]),
    .out1(in_reg_wire_7[137]),
    .out2(in_reg_wire_7[138]),
    .out3(in_reg_wire_7[139])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_35
  (
    .sel(conf_out[1823:1816]),
    .in0(in_reg_wire_6[35]),
    .in1(in_reg_wire_6[99]),
    .in2(in_reg_wire_6[163]),
    .in3(in_reg_wire_6[227]),
    .out0(in_reg_wire_7[140]),
    .out1(in_reg_wire_7[141]),
    .out2(in_reg_wire_7[142]),
    .out3(in_reg_wire_7[143])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_36
  (
    .sel(conf_out[1831:1824]),
    .in0(in_reg_wire_6[36]),
    .in1(in_reg_wire_6[100]),
    .in2(in_reg_wire_6[164]),
    .in3(in_reg_wire_6[228]),
    .out0(in_reg_wire_7[144]),
    .out1(in_reg_wire_7[145]),
    .out2(in_reg_wire_7[146]),
    .out3(in_reg_wire_7[147])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_37
  (
    .sel(conf_out[1839:1832]),
    .in0(in_reg_wire_6[37]),
    .in1(in_reg_wire_6[101]),
    .in2(in_reg_wire_6[165]),
    .in3(in_reg_wire_6[229]),
    .out0(in_reg_wire_7[148]),
    .out1(in_reg_wire_7[149]),
    .out2(in_reg_wire_7[150]),
    .out3(in_reg_wire_7[151])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_38
  (
    .sel(conf_out[1847:1840]),
    .in0(in_reg_wire_6[38]),
    .in1(in_reg_wire_6[102]),
    .in2(in_reg_wire_6[166]),
    .in3(in_reg_wire_6[230]),
    .out0(in_reg_wire_7[152]),
    .out1(in_reg_wire_7[153]),
    .out2(in_reg_wire_7[154]),
    .out3(in_reg_wire_7[155])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_39
  (
    .sel(conf_out[1855:1848]),
    .in0(in_reg_wire_6[39]),
    .in1(in_reg_wire_6[103]),
    .in2(in_reg_wire_6[167]),
    .in3(in_reg_wire_6[231]),
    .out0(in_reg_wire_7[156]),
    .out1(in_reg_wire_7[157]),
    .out2(in_reg_wire_7[158]),
    .out3(in_reg_wire_7[159])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_40
  (
    .sel(conf_out[1863:1856]),
    .in0(in_reg_wire_6[40]),
    .in1(in_reg_wire_6[104]),
    .in2(in_reg_wire_6[168]),
    .in3(in_reg_wire_6[232]),
    .out0(in_reg_wire_7[160]),
    .out1(in_reg_wire_7[161]),
    .out2(in_reg_wire_7[162]),
    .out3(in_reg_wire_7[163])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_41
  (
    .sel(conf_out[1871:1864]),
    .in0(in_reg_wire_6[41]),
    .in1(in_reg_wire_6[105]),
    .in2(in_reg_wire_6[169]),
    .in3(in_reg_wire_6[233]),
    .out0(in_reg_wire_7[164]),
    .out1(in_reg_wire_7[165]),
    .out2(in_reg_wire_7[166]),
    .out3(in_reg_wire_7[167])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_42
  (
    .sel(conf_out[1879:1872]),
    .in0(in_reg_wire_6[42]),
    .in1(in_reg_wire_6[106]),
    .in2(in_reg_wire_6[170]),
    .in3(in_reg_wire_6[234]),
    .out0(in_reg_wire_7[168]),
    .out1(in_reg_wire_7[169]),
    .out2(in_reg_wire_7[170]),
    .out3(in_reg_wire_7[171])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_43
  (
    .sel(conf_out[1887:1880]),
    .in0(in_reg_wire_6[43]),
    .in1(in_reg_wire_6[107]),
    .in2(in_reg_wire_6[171]),
    .in3(in_reg_wire_6[235]),
    .out0(in_reg_wire_7[172]),
    .out1(in_reg_wire_7[173]),
    .out2(in_reg_wire_7[174]),
    .out3(in_reg_wire_7[175])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_44
  (
    .sel(conf_out[1895:1888]),
    .in0(in_reg_wire_6[44]),
    .in1(in_reg_wire_6[108]),
    .in2(in_reg_wire_6[172]),
    .in3(in_reg_wire_6[236]),
    .out0(in_reg_wire_7[176]),
    .out1(in_reg_wire_7[177]),
    .out2(in_reg_wire_7[178]),
    .out3(in_reg_wire_7[179])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_45
  (
    .sel(conf_out[1903:1896]),
    .in0(in_reg_wire_6[45]),
    .in1(in_reg_wire_6[109]),
    .in2(in_reg_wire_6[173]),
    .in3(in_reg_wire_6[237]),
    .out0(in_reg_wire_7[180]),
    .out1(in_reg_wire_7[181]),
    .out2(in_reg_wire_7[182]),
    .out3(in_reg_wire_7[183])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_46
  (
    .sel(conf_out[1911:1904]),
    .in0(in_reg_wire_6[46]),
    .in1(in_reg_wire_6[110]),
    .in2(in_reg_wire_6[174]),
    .in3(in_reg_wire_6[238]),
    .out0(in_reg_wire_7[184]),
    .out1(in_reg_wire_7[185]),
    .out2(in_reg_wire_7[186]),
    .out3(in_reg_wire_7[187])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_47
  (
    .sel(conf_out[1919:1912]),
    .in0(in_reg_wire_6[47]),
    .in1(in_reg_wire_6[111]),
    .in2(in_reg_wire_6[175]),
    .in3(in_reg_wire_6[239]),
    .out0(in_reg_wire_7[188]),
    .out1(in_reg_wire_7[189]),
    .out2(in_reg_wire_7[190]),
    .out3(in_reg_wire_7[191])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_48
  (
    .sel(conf_out[1927:1920]),
    .in0(in_reg_wire_6[48]),
    .in1(in_reg_wire_6[112]),
    .in2(in_reg_wire_6[176]),
    .in3(in_reg_wire_6[240]),
    .out0(in_reg_wire_7[192]),
    .out1(in_reg_wire_7[193]),
    .out2(in_reg_wire_7[194]),
    .out3(in_reg_wire_7[195])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_49
  (
    .sel(conf_out[1935:1928]),
    .in0(in_reg_wire_6[49]),
    .in1(in_reg_wire_6[113]),
    .in2(in_reg_wire_6[177]),
    .in3(in_reg_wire_6[241]),
    .out0(in_reg_wire_7[196]),
    .out1(in_reg_wire_7[197]),
    .out2(in_reg_wire_7[198]),
    .out3(in_reg_wire_7[199])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_50
  (
    .sel(conf_out[1943:1936]),
    .in0(in_reg_wire_6[50]),
    .in1(in_reg_wire_6[114]),
    .in2(in_reg_wire_6[178]),
    .in3(in_reg_wire_6[242]),
    .out0(in_reg_wire_7[200]),
    .out1(in_reg_wire_7[201]),
    .out2(in_reg_wire_7[202]),
    .out3(in_reg_wire_7[203])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_51
  (
    .sel(conf_out[1951:1944]),
    .in0(in_reg_wire_6[51]),
    .in1(in_reg_wire_6[115]),
    .in2(in_reg_wire_6[179]),
    .in3(in_reg_wire_6[243]),
    .out0(in_reg_wire_7[204]),
    .out1(in_reg_wire_7[205]),
    .out2(in_reg_wire_7[206]),
    .out3(in_reg_wire_7[207])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_52
  (
    .sel(conf_out[1959:1952]),
    .in0(in_reg_wire_6[52]),
    .in1(in_reg_wire_6[116]),
    .in2(in_reg_wire_6[180]),
    .in3(in_reg_wire_6[244]),
    .out0(in_reg_wire_7[208]),
    .out1(in_reg_wire_7[209]),
    .out2(in_reg_wire_7[210]),
    .out3(in_reg_wire_7[211])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_53
  (
    .sel(conf_out[1967:1960]),
    .in0(in_reg_wire_6[53]),
    .in1(in_reg_wire_6[117]),
    .in2(in_reg_wire_6[181]),
    .in3(in_reg_wire_6[245]),
    .out0(in_reg_wire_7[212]),
    .out1(in_reg_wire_7[213]),
    .out2(in_reg_wire_7[214]),
    .out3(in_reg_wire_7[215])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_54
  (
    .sel(conf_out[1975:1968]),
    .in0(in_reg_wire_6[54]),
    .in1(in_reg_wire_6[118]),
    .in2(in_reg_wire_6[182]),
    .in3(in_reg_wire_6[246]),
    .out0(in_reg_wire_7[216]),
    .out1(in_reg_wire_7[217]),
    .out2(in_reg_wire_7[218]),
    .out3(in_reg_wire_7[219])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_55
  (
    .sel(conf_out[1983:1976]),
    .in0(in_reg_wire_6[55]),
    .in1(in_reg_wire_6[119]),
    .in2(in_reg_wire_6[183]),
    .in3(in_reg_wire_6[247]),
    .out0(in_reg_wire_7[220]),
    .out1(in_reg_wire_7[221]),
    .out2(in_reg_wire_7[222]),
    .out3(in_reg_wire_7[223])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_56
  (
    .sel(conf_out[1991:1984]),
    .in0(in_reg_wire_6[56]),
    .in1(in_reg_wire_6[120]),
    .in2(in_reg_wire_6[184]),
    .in3(in_reg_wire_6[248]),
    .out0(in_reg_wire_7[224]),
    .out1(in_reg_wire_7[225]),
    .out2(in_reg_wire_7[226]),
    .out3(in_reg_wire_7[227])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_57
  (
    .sel(conf_out[1999:1992]),
    .in0(in_reg_wire_6[57]),
    .in1(in_reg_wire_6[121]),
    .in2(in_reg_wire_6[185]),
    .in3(in_reg_wire_6[249]),
    .out0(in_reg_wire_7[228]),
    .out1(in_reg_wire_7[229]),
    .out2(in_reg_wire_7[230]),
    .out3(in_reg_wire_7[231])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_58
  (
    .sel(conf_out[2007:2000]),
    .in0(in_reg_wire_6[58]),
    .in1(in_reg_wire_6[122]),
    .in2(in_reg_wire_6[186]),
    .in3(in_reg_wire_6[250]),
    .out0(in_reg_wire_7[232]),
    .out1(in_reg_wire_7[233]),
    .out2(in_reg_wire_7[234]),
    .out3(in_reg_wire_7[235])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_59
  (
    .sel(conf_out[2015:2008]),
    .in0(in_reg_wire_6[59]),
    .in1(in_reg_wire_6[123]),
    .in2(in_reg_wire_6[187]),
    .in3(in_reg_wire_6[251]),
    .out0(in_reg_wire_7[236]),
    .out1(in_reg_wire_7[237]),
    .out2(in_reg_wire_7[238]),
    .out3(in_reg_wire_7[239])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_60
  (
    .sel(conf_out[2023:2016]),
    .in0(in_reg_wire_6[60]),
    .in1(in_reg_wire_6[124]),
    .in2(in_reg_wire_6[188]),
    .in3(in_reg_wire_6[252]),
    .out0(in_reg_wire_7[240]),
    .out1(in_reg_wire_7[241]),
    .out2(in_reg_wire_7[242]),
    .out3(in_reg_wire_7[243])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_61
  (
    .sel(conf_out[2031:2024]),
    .in0(in_reg_wire_6[61]),
    .in1(in_reg_wire_6[125]),
    .in2(in_reg_wire_6[189]),
    .in3(in_reg_wire_6[253]),
    .out0(in_reg_wire_7[244]),
    .out1(in_reg_wire_7[245]),
    .out2(in_reg_wire_7[246]),
    .out3(in_reg_wire_7[247])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_62
  (
    .sel(conf_out[2039:2032]),
    .in0(in_reg_wire_6[62]),
    .in1(in_reg_wire_6[126]),
    .in2(in_reg_wire_6[190]),
    .in3(in_reg_wire_6[254]),
    .out0(in_reg_wire_7[248]),
    .out1(in_reg_wire_7[249]),
    .out2(in_reg_wire_7[250]),
    .out3(in_reg_wire_7[251])
  );


  switch_box4x4
  #(
    .WIDTH(WIDTH)
  )
  sw_3_63
  (
    .sel(conf_out[2047:2040]),
    .in0(in_reg_wire_6[63]),
    .in1(in_reg_wire_6[127]),
    .in2(in_reg_wire_6[191]),
    .in3(in_reg_wire_6[255]),
    .out0(in_reg_wire_7[252]),
    .out1(in_reg_wire_7[253]),
    .out2(in_reg_wire_7[254]),
    .out3(in_reg_wire_7[255])
  );

endmodule