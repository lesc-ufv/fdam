module reg_tree_4_66_2 #
(
  parameter DATA_WIDTH = 16
)
(
  input clk,
  input [DATA_WIDTH-1:0] in,
  output [DATA_WIDTH-1:0] out_0,
  output [DATA_WIDTH-1:0] out_1,
  output [DATA_WIDTH-1:0] out_2,
  output [DATA_WIDTH-1:0] out_3,
  output [DATA_WIDTH-1:0] out_4,
  output [DATA_WIDTH-1:0] out_5,
  output [DATA_WIDTH-1:0] out_6,
  output [DATA_WIDTH-1:0] out_7,
  output [DATA_WIDTH-1:0] out_8,
  output [DATA_WIDTH-1:0] out_9,
  output [DATA_WIDTH-1:0] out_10,
  output [DATA_WIDTH-1:0] out_11,
  output [DATA_WIDTH-1:0] out_12,
  output [DATA_WIDTH-1:0] out_13,
  output [DATA_WIDTH-1:0] out_14,
  output [DATA_WIDTH-1:0] out_15,
  output [DATA_WIDTH-1:0] out_16,
  output [DATA_WIDTH-1:0] out_17,
  output [DATA_WIDTH-1:0] out_18,
  output [DATA_WIDTH-1:0] out_19,
  output [DATA_WIDTH-1:0] out_20,
  output [DATA_WIDTH-1:0] out_21,
  output [DATA_WIDTH-1:0] out_22,
  output [DATA_WIDTH-1:0] out_23,
  output [DATA_WIDTH-1:0] out_24,
  output [DATA_WIDTH-1:0] out_25,
  output [DATA_WIDTH-1:0] out_26,
  output [DATA_WIDTH-1:0] out_27,
  output [DATA_WIDTH-1:0] out_28,
  output [DATA_WIDTH-1:0] out_29,
  output [DATA_WIDTH-1:0] out_30,
  output [DATA_WIDTH-1:0] out_31,
  output [DATA_WIDTH-1:0] out_32,
  output [DATA_WIDTH-1:0] out_33,
  output [DATA_WIDTH-1:0] out_34,
  output [DATA_WIDTH-1:0] out_35,
  output [DATA_WIDTH-1:0] out_36,
  output [DATA_WIDTH-1:0] out_37,
  output [DATA_WIDTH-1:0] out_38,
  output [DATA_WIDTH-1:0] out_39,
  output [DATA_WIDTH-1:0] out_40,
  output [DATA_WIDTH-1:0] out_41,
  output [DATA_WIDTH-1:0] out_42,
  output [DATA_WIDTH-1:0] out_43,
  output [DATA_WIDTH-1:0] out_44,
  output [DATA_WIDTH-1:0] out_45,
  output [DATA_WIDTH-1:0] out_46,
  output [DATA_WIDTH-1:0] out_47,
  output [DATA_WIDTH-1:0] out_48,
  output [DATA_WIDTH-1:0] out_49,
  output [DATA_WIDTH-1:0] out_50,
  output [DATA_WIDTH-1:0] out_51,
  output [DATA_WIDTH-1:0] out_52,
  output [DATA_WIDTH-1:0] out_53,
  output [DATA_WIDTH-1:0] out_54,
  output [DATA_WIDTH-1:0] out_55,
  output [DATA_WIDTH-1:0] out_56,
  output [DATA_WIDTH-1:0] out_57,
  output [DATA_WIDTH-1:0] out_58,
  output [DATA_WIDTH-1:0] out_59,
  output [DATA_WIDTH-1:0] out_60,
  output [DATA_WIDTH-1:0] out_61,
  output [DATA_WIDTH-1:0] out_62,
  output [DATA_WIDTH-1:0] out_63,
  output [DATA_WIDTH-1:0] out_64,
  output [DATA_WIDTH-1:0] out_65
);

  reg [DATA_WIDTH-1:0] r0;
  reg [DATA_WIDTH-1:0] r1;
  reg [DATA_WIDTH-1:0] r2;
  reg [DATA_WIDTH-1:0] r3;
  reg [DATA_WIDTH-1:0] r4;
  reg [DATA_WIDTH-1:0] r5;
  reg [DATA_WIDTH-1:0] r6;
  reg [DATA_WIDTH-1:0] r7;
  reg [DATA_WIDTH-1:0] r8;
  reg [DATA_WIDTH-1:0] r9;
  reg [DATA_WIDTH-1:0] r10;
  reg [DATA_WIDTH-1:0] r11;
  reg [DATA_WIDTH-1:0] r12;
  reg [DATA_WIDTH-1:0] r13;
  reg [DATA_WIDTH-1:0] r14;
  reg [DATA_WIDTH-1:0] r15;
  reg [DATA_WIDTH-1:0] r16;
  reg [DATA_WIDTH-1:0] r17;
  reg [DATA_WIDTH-1:0] r18;
  reg [DATA_WIDTH-1:0] r19;
  reg [DATA_WIDTH-1:0] r20;
  reg [DATA_WIDTH-1:0] r21;
  reg [DATA_WIDTH-1:0] r22;
  reg [DATA_WIDTH-1:0] r23;
  reg [DATA_WIDTH-1:0] r24;
  reg [DATA_WIDTH-1:0] r25;
  reg [DATA_WIDTH-1:0] r26;
  reg [DATA_WIDTH-1:0] r27;
  reg [DATA_WIDTH-1:0] r28;
  reg [DATA_WIDTH-1:0] r29;
  reg [DATA_WIDTH-1:0] r30;
  reg [DATA_WIDTH-1:0] r31;
  reg [DATA_WIDTH-1:0] r32;
  reg [DATA_WIDTH-1:0] r33;
  reg [DATA_WIDTH-1:0] r34;
  reg [DATA_WIDTH-1:0] r35;
  reg [DATA_WIDTH-1:0] r36;
  reg [DATA_WIDTH-1:0] r37;
  reg [DATA_WIDTH-1:0] r38;
  reg [DATA_WIDTH-1:0] r39;
  reg [DATA_WIDTH-1:0] r40;
  reg [DATA_WIDTH-1:0] r41;
  reg [DATA_WIDTH-1:0] r42;
  reg [DATA_WIDTH-1:0] r43;
  reg [DATA_WIDTH-1:0] r44;
  reg [DATA_WIDTH-1:0] r45;
  reg [DATA_WIDTH-1:0] r46;
  reg [DATA_WIDTH-1:0] r47;
  reg [DATA_WIDTH-1:0] r48;
  reg [DATA_WIDTH-1:0] r49;
  reg [DATA_WIDTH-1:0] r50;
  reg [DATA_WIDTH-1:0] r51;
  reg [DATA_WIDTH-1:0] r52;
  reg [DATA_WIDTH-1:0] r53;
  reg [DATA_WIDTH-1:0] r54;
  reg [DATA_WIDTH-1:0] r55;
  reg [DATA_WIDTH-1:0] r56;
  reg [DATA_WIDTH-1:0] r57;
  reg [DATA_WIDTH-1:0] r58;
  reg [DATA_WIDTH-1:0] r59;
  reg [DATA_WIDTH-1:0] r60;
  reg [DATA_WIDTH-1:0] r61;
  reg [DATA_WIDTH-1:0] r62;
  reg [DATA_WIDTH-1:0] r63;
  reg [DATA_WIDTH-1:0] r64;
  reg [DATA_WIDTH-1:0] r65;
  reg [DATA_WIDTH-1:0] r66;
  reg [DATA_WIDTH-1:0] r67;
  reg [DATA_WIDTH-1:0] r68;
  reg [DATA_WIDTH-1:0] r69;
  reg [DATA_WIDTH-1:0] r70;
  reg [DATA_WIDTH-1:0] r71;
  reg [DATA_WIDTH-1:0] r72;
  reg [DATA_WIDTH-1:0] r73;
  reg [DATA_WIDTH-1:0] r74;
  reg [DATA_WIDTH-1:0] r75;
  reg [DATA_WIDTH-1:0] r76;
  reg [DATA_WIDTH-1:0] r77;
  reg [DATA_WIDTH-1:0] r78;
  reg [DATA_WIDTH-1:0] r79;
  reg [DATA_WIDTH-1:0] r80;
  reg [DATA_WIDTH-1:0] r81;
  reg [DATA_WIDTH-1:0] r82;
  reg [DATA_WIDTH-1:0] r83;
  reg [DATA_WIDTH-1:0] r84;
  reg [DATA_WIDTH-1:0] r85;
  reg [DATA_WIDTH-1:0] r86;
  reg [DATA_WIDTH-1:0] r87;
  reg [DATA_WIDTH-1:0] r88;
  reg [DATA_WIDTH-1:0] r89;
  reg [DATA_WIDTH-1:0] r90;
  reg [DATA_WIDTH-1:0] r91;
  reg [DATA_WIDTH-1:0] r92;
  reg [DATA_WIDTH-1:0] r93;
  reg [DATA_WIDTH-1:0] r94;
  reg [DATA_WIDTH-1:0] r95;
  reg [DATA_WIDTH-1:0] r96;
  reg [DATA_WIDTH-1:0] r97;
  reg [DATA_WIDTH-1:0] r98;
  reg [DATA_WIDTH-1:0] r99;
  reg [DATA_WIDTH-1:0] r100;
  reg [DATA_WIDTH-1:0] r101;
  reg [DATA_WIDTH-1:0] r102;
  reg [DATA_WIDTH-1:0] r103;
  reg [DATA_WIDTH-1:0] r104;
  reg [DATA_WIDTH-1:0] r105;
  reg [DATA_WIDTH-1:0] r106;
  reg [DATA_WIDTH-1:0] r107;
  reg [DATA_WIDTH-1:0] r108;
  reg [DATA_WIDTH-1:0] r109;
  reg [DATA_WIDTH-1:0] r110;
  reg [DATA_WIDTH-1:0] r111;
  reg [DATA_WIDTH-1:0] r112;
  reg [DATA_WIDTH-1:0] r113;
  reg [DATA_WIDTH-1:0] r114;
  reg [DATA_WIDTH-1:0] r115;
  reg [DATA_WIDTH-1:0] r116;
  reg [DATA_WIDTH-1:0] r117;
  reg [DATA_WIDTH-1:0] r118;
  reg [DATA_WIDTH-1:0] r119;
  reg [DATA_WIDTH-1:0] r120;
  reg [DATA_WIDTH-1:0] r121;
  reg [DATA_WIDTH-1:0] r122;
  reg [DATA_WIDTH-1:0] r123;
  reg [DATA_WIDTH-1:0] r124;
  reg [DATA_WIDTH-1:0] r125;
  reg [DATA_WIDTH-1:0] r126;
  reg [DATA_WIDTH-1:0] r127;
  reg [DATA_WIDTH-1:0] r128;
  reg [DATA_WIDTH-1:0] r129;
  reg [DATA_WIDTH-1:0] r130;
  reg [DATA_WIDTH-1:0] r131;
  reg [DATA_WIDTH-1:0] r132;
  reg [DATA_WIDTH-1:0] r133;
  reg [DATA_WIDTH-1:0] r134;
  reg [DATA_WIDTH-1:0] r135;
  reg [DATA_WIDTH-1:0] r136;
  reg [DATA_WIDTH-1:0] r137;
  reg [DATA_WIDTH-1:0] r138;
  reg [DATA_WIDTH-1:0] r139;
  reg [DATA_WIDTH-1:0] r140;
  reg [DATA_WIDTH-1:0] r141;
  reg [DATA_WIDTH-1:0] r142;
  reg [DATA_WIDTH-1:0] r143;
  reg [DATA_WIDTH-1:0] r144;
  reg [DATA_WIDTH-1:0] r145;
  reg [DATA_WIDTH-1:0] r146;
  reg [DATA_WIDTH-1:0] r147;
  reg [DATA_WIDTH-1:0] r148;
  reg [DATA_WIDTH-1:0] r149;
  reg [DATA_WIDTH-1:0] r150;
  reg [DATA_WIDTH-1:0] r151;
  reg [DATA_WIDTH-1:0] r152;
  reg [DATA_WIDTH-1:0] r153;
  reg [DATA_WIDTH-1:0] r154;
  reg [DATA_WIDTH-1:0] r155;
  reg [DATA_WIDTH-1:0] r156;
  reg [DATA_WIDTH-1:0] r157;
  reg [DATA_WIDTH-1:0] r158;
  reg [DATA_WIDTH-1:0] r159;
  reg [DATA_WIDTH-1:0] r160;
  reg [DATA_WIDTH-1:0] r161;
  reg [DATA_WIDTH-1:0] r162;
  reg [DATA_WIDTH-1:0] r163;
  reg [DATA_WIDTH-1:0] r164;
  reg [DATA_WIDTH-1:0] r165;
  reg [DATA_WIDTH-1:0] r166;
  reg [DATA_WIDTH-1:0] r167;
  reg [DATA_WIDTH-1:0] r168;
  reg [DATA_WIDTH-1:0] r169;
  reg [DATA_WIDTH-1:0] r170;
  reg [DATA_WIDTH-1:0] r171;
  reg [DATA_WIDTH-1:0] r172;
  reg [DATA_WIDTH-1:0] r173;
  reg [DATA_WIDTH-1:0] r174;
  reg [DATA_WIDTH-1:0] r175;
  reg [DATA_WIDTH-1:0] r176;
  reg [DATA_WIDTH-1:0] r177;
  reg [DATA_WIDTH-1:0] r178;
  reg [DATA_WIDTH-1:0] r179;
  reg [DATA_WIDTH-1:0] r180;
  reg [DATA_WIDTH-1:0] r181;
  reg [DATA_WIDTH-1:0] r182;
  reg [DATA_WIDTH-1:0] r183;
  reg [DATA_WIDTH-1:0] r184;
  reg [DATA_WIDTH-1:0] r185;
  reg [DATA_WIDTH-1:0] r186;
  reg [DATA_WIDTH-1:0] r187;
  reg [DATA_WIDTH-1:0] r188;
  reg [DATA_WIDTH-1:0] r189;
  reg [DATA_WIDTH-1:0] r190;
  reg [DATA_WIDTH-1:0] r191;
  reg [DATA_WIDTH-1:0] r192;
  reg [DATA_WIDTH-1:0] r193;
  reg [DATA_WIDTH-1:0] r194;
  reg [DATA_WIDTH-1:0] r195;
  reg [DATA_WIDTH-1:0] r196;
  reg [DATA_WIDTH-1:0] r197;
  reg [DATA_WIDTH-1:0] r198;
  reg [DATA_WIDTH-1:0] r199;
  reg [DATA_WIDTH-1:0] r200;
  reg [DATA_WIDTH-1:0] r201;
  reg [DATA_WIDTH-1:0] r202;
  reg [DATA_WIDTH-1:0] r203;
  reg [DATA_WIDTH-1:0] r204;
  reg [DATA_WIDTH-1:0] r205;
  reg [DATA_WIDTH-1:0] r206;
  reg [DATA_WIDTH-1:0] r207;
  reg [DATA_WIDTH-1:0] r208;
  reg [DATA_WIDTH-1:0] r209;
  reg [DATA_WIDTH-1:0] r210;
  reg [DATA_WIDTH-1:0] r211;
  reg [DATA_WIDTH-1:0] r212;
  reg [DATA_WIDTH-1:0] r213;
  reg [DATA_WIDTH-1:0] r214;
  reg [DATA_WIDTH-1:0] r215;
  reg [DATA_WIDTH-1:0] r216;
  reg [DATA_WIDTH-1:0] r217;
  reg [DATA_WIDTH-1:0] r218;
  reg [DATA_WIDTH-1:0] r219;
  reg [DATA_WIDTH-1:0] r220;
  reg [DATA_WIDTH-1:0] r221;
  reg [DATA_WIDTH-1:0] r222;

  initial begin
    r0 = 0;
    r1 = 0;
    r2 = 0;
    r3 = 0;
    r4 = 0;
    r5 = 0;
    r6 = 0;
    r7 = 0;
    r8 = 0;
    r9 = 0;
    r10 = 0;
    r11 = 0;
    r12 = 0;
    r13 = 0;
    r14 = 0;
    r15 = 0;
    r16 = 0;
    r17 = 0;
    r18 = 0;
    r19 = 0;
    r20 = 0;
    r21 = 0;
    r22 = 0;
    r23 = 0;
    r24 = 0;
    r25 = 0;
    r26 = 0;
    r27 = 0;
    r28 = 0;
    r29 = 0;
    r30 = 0;
    r31 = 0;
    r32 = 0;
    r33 = 0;
    r34 = 0;
    r35 = 0;
    r36 = 0;
    r37 = 0;
    r38 = 0;
    r39 = 0;
    r40 = 0;
    r41 = 0;
    r42 = 0;
    r43 = 0;
    r44 = 0;
    r45 = 0;
    r46 = 0;
    r47 = 0;
    r48 = 0;
    r49 = 0;
    r50 = 0;
    r51 = 0;
    r52 = 0;
    r53 = 0;
    r54 = 0;
    r55 = 0;
    r56 = 0;
    r57 = 0;
    r58 = 0;
    r59 = 0;
    r60 = 0;
    r61 = 0;
    r62 = 0;
    r63 = 0;
    r64 = 0;
    r65 = 0;
    r66 = 0;
    r67 = 0;
    r68 = 0;
    r69 = 0;
    r70 = 0;
    r71 = 0;
    r72 = 0;
    r73 = 0;
    r74 = 0;
    r75 = 0;
    r76 = 0;
    r77 = 0;
    r78 = 0;
    r79 = 0;
    r80 = 0;
    r81 = 0;
    r82 = 0;
    r83 = 0;
    r84 = 0;
    r85 = 0;
    r86 = 0;
    r87 = 0;
    r88 = 0;
    r89 = 0;
    r90 = 0;
    r91 = 0;
    r92 = 0;
    r93 = 0;
    r94 = 0;
    r95 = 0;
    r96 = 0;
    r97 = 0;
    r98 = 0;
    r99 = 0;
    r100 = 0;
    r101 = 0;
    r102 = 0;
    r103 = 0;
    r104 = 0;
    r105 = 0;
    r106 = 0;
    r107 = 0;
    r108 = 0;
    r109 = 0;
    r110 = 0;
    r111 = 0;
    r112 = 0;
    r113 = 0;
    r114 = 0;
    r115 = 0;
    r116 = 0;
    r117 = 0;
    r118 = 0;
    r119 = 0;
    r120 = 0;
    r121 = 0;
    r122 = 0;
    r123 = 0;
    r124 = 0;
    r125 = 0;
    r126 = 0;
    r127 = 0;
    r128 = 0;
    r129 = 0;
    r130 = 0;
    r131 = 0;
    r132 = 0;
    r133 = 0;
    r134 = 0;
    r135 = 0;
    r136 = 0;
    r137 = 0;
    r138 = 0;
    r139 = 0;
    r140 = 0;
    r141 = 0;
    r142 = 0;
    r143 = 0;
    r144 = 0;
    r145 = 0;
    r146 = 0;
    r147 = 0;
    r148 = 0;
    r149 = 0;
    r150 = 0;
    r151 = 0;
    r152 = 0;
    r153 = 0;
    r154 = 0;
    r155 = 0;
    r156 = 0;
    r157 = 0;
    r158 = 0;
    r159 = 0;
    r160 = 0;
    r161 = 0;
    r162 = 0;
    r163 = 0;
    r164 = 0;
    r165 = 0;
    r166 = 0;
    r167 = 0;
    r168 = 0;
    r169 = 0;
    r170 = 0;
    r171 = 0;
    r172 = 0;
    r173 = 0;
    r174 = 0;
    r175 = 0;
    r176 = 0;
    r177 = 0;
    r178 = 0;
    r179 = 0;
    r180 = 0;
    r181 = 0;
    r182 = 0;
    r183 = 0;
    r184 = 0;
    r185 = 0;
    r186 = 0;
    r187 = 0;
    r188 = 0;
    r189 = 0;
    r190 = 0;
    r191 = 0;
    r192 = 0;
    r193 = 0;
    r194 = 0;
    r195 = 0;
    r196 = 0;
    r197 = 0;
    r198 = 0;
    r199 = 0;
    r200 = 0;
    r201 = 0;
    r202 = 0;
    r203 = 0;
    r204 = 0;
    r205 = 0;
    r206 = 0;
    r207 = 0;
    r208 = 0;
    r209 = 0;
    r210 = 0;
    r211 = 0;
    r212 = 0;
    r213 = 0;
    r214 = 0;
    r215 = 0;
    r216 = 0;
    r217 = 0;
    r218 = 0;
    r219 = 0;
    r220 = 0;
    r221 = 0;
    r222 = 0;

  end



  always @(posedge clk) begin
    r0 <= in;
    r1 <= r0;
    r2 <= r0;
    r3 <= r1;
    r4 <= r1;
    r5 <= r1;
    r6 <= r1;
    r7 <= r2;
    r8 <= r3;
    r9 <= r3;
    r10 <= r3;
    r11 <= r3;
    r12 <= r4;
    r13 <= r4;
    r14 <= r4;
    r15 <= r4;
    r16 <= r5;
    r17 <= r5;
    r18 <= r5;
    r19 <= r5;
    r20 <= r6;
    r21 <= r6;
    r22 <= r6;
    r23 <= r6;
    r24 <= r7;
    r25 <= r8;
    r26 <= r8;
    r27 <= r8;
    r28 <= r8;
    r29 <= r9;
    r30 <= r9;
    r31 <= r9;
    r32 <= r9;
    r33 <= r10;
    r34 <= r10;
    r35 <= r10;
    r36 <= r10;
    r37 <= r11;
    r38 <= r11;
    r39 <= r11;
    r40 <= r11;
    r41 <= r12;
    r42 <= r12;
    r43 <= r12;
    r44 <= r12;
    r45 <= r13;
    r46 <= r13;
    r47 <= r13;
    r48 <= r13;
    r49 <= r14;
    r50 <= r14;
    r51 <= r14;
    r52 <= r14;
    r53 <= r15;
    r54 <= r15;
    r55 <= r15;
    r56 <= r15;
    r57 <= r16;
    r58 <= r16;
    r59 <= r16;
    r60 <= r16;
    r61 <= r17;
    r62 <= r17;
    r63 <= r17;
    r64 <= r17;
    r65 <= r18;
    r66 <= r18;
    r67 <= r18;
    r68 <= r18;
    r69 <= r19;
    r70 <= r19;
    r71 <= r19;
    r72 <= r19;
    r73 <= r20;
    r74 <= r20;
    r75 <= r20;
    r76 <= r20;
    r77 <= r21;
    r78 <= r21;
    r79 <= r21;
    r80 <= r21;
    r81 <= r22;
    r82 <= r22;
    r83 <= r22;
    r84 <= r22;
    r85 <= r23;
    r86 <= r23;
    r87 <= r23;
    r88 <= r23;
    r89 <= r24;
    r90 <= r24;
    r91 <= r25;
    r92 <= r26;
    r93 <= r27;
    r94 <= r28;
    r95 <= r29;
    r96 <= r30;
    r97 <= r31;
    r98 <= r32;
    r99 <= r33;
    r100 <= r34;
    r101 <= r35;
    r102 <= r36;
    r103 <= r37;
    r104 <= r38;
    r105 <= r39;
    r106 <= r40;
    r107 <= r41;
    r108 <= r42;
    r109 <= r43;
    r110 <= r44;
    r111 <= r45;
    r112 <= r46;
    r113 <= r47;
    r114 <= r48;
    r115 <= r49;
    r116 <= r50;
    r117 <= r51;
    r118 <= r52;
    r119 <= r53;
    r120 <= r54;
    r121 <= r55;
    r122 <= r56;
    r123 <= r57;
    r124 <= r58;
    r125 <= r59;
    r126 <= r60;
    r127 <= r61;
    r128 <= r62;
    r129 <= r63;
    r130 <= r64;
    r131 <= r65;
    r132 <= r66;
    r133 <= r67;
    r134 <= r68;
    r135 <= r69;
    r136 <= r70;
    r137 <= r71;
    r138 <= r72;
    r139 <= r73;
    r140 <= r74;
    r141 <= r75;
    r142 <= r76;
    r143 <= r77;
    r144 <= r78;
    r145 <= r79;
    r146 <= r80;
    r147 <= r81;
    r148 <= r82;
    r149 <= r83;
    r150 <= r84;
    r151 <= r85;
    r152 <= r86;
    r153 <= r87;
    r154 <= r88;
    r155 <= r89;
    r156 <= r90;
    r157 <= r91;
    r158 <= r92;
    r159 <= r93;
    r160 <= r94;
    r161 <= r95;
    r162 <= r96;
    r163 <= r97;
    r164 <= r98;
    r165 <= r99;
    r166 <= r100;
    r167 <= r101;
    r168 <= r102;
    r169 <= r103;
    r170 <= r104;
    r171 <= r105;
    r172 <= r106;
    r173 <= r107;
    r174 <= r108;
    r175 <= r109;
    r176 <= r110;
    r177 <= r111;
    r178 <= r112;
    r179 <= r113;
    r180 <= r114;
    r181 <= r115;
    r182 <= r116;
    r183 <= r117;
    r184 <= r118;
    r185 <= r119;
    r186 <= r120;
    r187 <= r121;
    r188 <= r122;
    r189 <= r123;
    r190 <= r124;
    r191 <= r125;
    r192 <= r126;
    r193 <= r127;
    r194 <= r128;
    r195 <= r129;
    r196 <= r130;
    r197 <= r131;
    r198 <= r132;
    r199 <= r133;
    r200 <= r134;
    r201 <= r135;
    r202 <= r136;
    r203 <= r137;
    r204 <= r138;
    r205 <= r139;
    r206 <= r140;
    r207 <= r141;
    r208 <= r142;
    r209 <= r143;
    r210 <= r144;
    r211 <= r145;
    r212 <= r146;
    r213 <= r147;
    r214 <= r148;
    r215 <= r149;
    r216 <= r150;
    r217 <= r151;
    r218 <= r152;
    r219 <= r153;
    r220 <= r154;
    r221 <= r155;
    r222 <= r156;

  end

  assign out_0 = r157;
  assign out_1 = r158;
  assign out_2 = r159;
  assign out_3 = r160;
  assign out_4 = r161;
  assign out_5 = r162;
  assign out_6 = r163;
  assign out_7 = r164;
  assign out_8 = r165;
  assign out_9 = r166;
  assign out_10 = r167;
  assign out_11 = r168;
  assign out_12 = r169;
  assign out_13 = r170;
  assign out_14 = r171;
  assign out_15 = r172;
  assign out_16 = r173;
  assign out_17 = r174;
  assign out_18 = r175;
  assign out_19 = r176;
  assign out_20 = r177;
  assign out_21 = r178;
  assign out_22 = r179;
  assign out_23 = r180;
  assign out_24 = r181;
  assign out_25 = r182;
  assign out_26 = r183;
  assign out_27 = r184;
  assign out_28 = r185;
  assign out_29 = r186;
  assign out_30 = r187;
  assign out_31 = r188;
  assign out_32 = r189;
  assign out_33 = r190;
  assign out_34 = r191;
  assign out_35 = r192;
  assign out_36 = r193;
  assign out_37 = r194;
  assign out_38 = r195;
  assign out_39 = r196;
  assign out_40 = r197;
  assign out_41 = r198;
  assign out_42 = r199;
  assign out_43 = r200;
  assign out_44 = r201;
  assign out_45 = r202;
  assign out_46 = r203;
  assign out_47 = r204;
  assign out_48 = r205;
  assign out_49 = r206;
  assign out_50 = r207;
  assign out_51 = r208;
  assign out_52 = r209;
  assign out_53 = r210;
  assign out_54 = r211;
  assign out_55 = r212;
  assign out_56 = r213;
  assign out_57 = r214;
  assign out_58 = r215;
  assign out_59 = r216;
  assign out_60 = r217;
  assign out_61 = r218;
  assign out_62 = r219;
  assign out_63 = r220;
  assign out_64 = r221;
  assign out_65 = r222;

endmodule